// niosII_system.v

// Generated using ACDS version 12.1sp1 243 at 2017.02.19.16:32:03

`timescale 1 ps / 1 ps
module niosII_system (
		input  wire        audio_core_external_interface_ADCDAT,                                  //          audio_core_external_interface.ADCDAT
		input  wire        audio_core_external_interface_ADCLRCK,                                 //                                       .ADCLRCK
		input  wire        audio_core_external_interface_BCLK,                                    //                                       .BCLK
		output wire        audio_core_external_interface_DACDAT,                                  //                                       .DACDAT
		input  wire        audio_core_external_interface_DACLRCK,                                 //                                       .DACLRCK
		input  wire        cancel_button_external_connection_export,                              //      cancel_button_external_connection.export
		inout  wire        audio_config_external_interface_SDAT,                                  //        audio_config_external_interface.SDAT
		output wire        audio_config_external_interface_SCLK,                                  //                                       .SCLK
		input  wire        clock_27mhz_clk_in_clk,                                                //                     clock_27mhz_clk_in.clk
		output wire [7:0]  red_leds_external_connection_export,                                   //           red_leds_external_connection.export
		input  wire        remove_button_external_connection_export,                              //      remove_button_external_connection.export
		input  wire        switch_external_connection_export,                                     //             switch_external_connection.export
		input  wire        clk_clk,                                                               //                                    clk.clk
		output wire [7:0]  green_leds_external_connection_export,                                 //         green_leds_external_connection.export
		inout  wire [15:0] sram_external_interface_DQ,                                            //                sram_external_interface.DQ
		output wire [17:0] sram_external_interface_ADDR,                                          //                                       .ADDR
		output wire        sram_external_interface_LB_N,                                          //                                       .LB_N
		output wire        sram_external_interface_UB_N,                                          //                                       .UB_N
		output wire        sram_external_interface_CE_N,                                          //                                       .CE_N
		output wire        sram_external_interface_OE_N,                                          //                                       .OE_N
		output wire        sram_external_interface_WE_N,                                          //                                       .WE_N
		inout  wire        barcode_scanner_ps2_external_interface_CLK,                            // barcode_scanner_ps2_external_interface.CLK
		inout  wire        barcode_scanner_ps2_external_interface_DAT,                            //                                       .DAT
		output wire [11:0] sdram_wire_addr,                                                       //                             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                                         //                                       .ba
		output wire        sdram_wire_cas_n,                                                      //                                       .cas_n
		output wire        sdram_wire_cke,                                                        //                                       .cke
		output wire        sdram_wire_cs_n,                                                       //                                       .cs_n
		inout  wire [15:0] sdram_wire_dq,                                                         //                                       .dq
		output wire [1:0]  sdram_wire_dqm,                                                        //                                       .dqm
		output wire        sdram_wire_ras_n,                                                      //                                       .ras_n
		output wire        sdram_wire_we_n,                                                       //                                       .we_n
		output wire        main_pll_sdram_clk_clk,                                                //                     main_pll_sdram_clk.clk
		input  wire        reset_reset_n,                                                         //                                  reset.reset_n
		inout  wire [15:0] dm9000a_if_ethernet_s1_export_DATA,                                    //          dm9000a_if_ethernet_s1_export.DATA
		output wire        dm9000a_if_ethernet_s1_export_CMD,                                     //                                       .CMD
		output wire        dm9000a_if_ethernet_s1_export_RD_N,                                    //                                       .RD_N
		output wire        dm9000a_if_ethernet_s1_export_WR_N,                                    //                                       .WR_N
		output wire        dm9000a_if_ethernet_s1_export_CS_N,                                    //                                       .CS_N
		output wire        dm9000a_if_ethernet_s1_export_RST_N,                                   //                                       .RST_N
		input  wire        dm9000a_if_ethernet_s1_export_INT,                                     //                                       .INT
		output wire        dm9000a_if_ethernet_s1_export_CLK,                                     //                                       .CLK
		inout  wire [7:0]  character_lcd_external_interface_DATA,                                 //       character_lcd_external_interface.DATA
		output wire        character_lcd_external_interface_ON,                                   //                                       .ON
		output wire        character_lcd_external_interface_BLON,                                 //                                       .BLON
		output wire        character_lcd_external_interface_EN,                                   //                                       .EN
		output wire        character_lcd_external_interface_RS,                                   //                                       .RS
		output wire        character_lcd_external_interface_RW,                                   //                                       .RW
		input  wire        add_button_external_connection_export,                                 //         add_button_external_connection.export
		output wire [0:0]  tristate_conduit_bridge_out_tristate_controller_tcm_read_n_out,        //            tristate_conduit_bridge_out.tristate_controller_tcm_read_n_out
		output wire [21:0] tristate_conduit_bridge_out_tristate_controller_tcm_address_out,       //                                       .tristate_controller_tcm_address_out
		inout  wire [7:0]  tristate_conduit_bridge_out_tristate_controller_tcm_data_out,          //                                       .tristate_controller_tcm_data_out
		output wire [0:0]  tristate_conduit_bridge_out_tristate_controller_tcm_byteenable_out,    //                                       .tristate_controller_tcm_byteenable_out
		output wire [0:0]  tristate_conduit_bridge_out_tristate_controller_tcm_begintransfer_out, //                                       .tristate_controller_tcm_begintransfer_out
		output wire [0:0]  tristate_conduit_bridge_out_tristate_controller_tcm_write_n_out,       //                                       .tristate_controller_tcm_write_n_out
		output wire [0:0]  tristate_conduit_bridge_out_tristate_controller_tcm_chipselect_n_out,  //                                       .tristate_controller_tcm_chipselect_n_out
		input  wire        clock_27mhz_clk_in_reset_reset_n                                       //               clock_27mhz_clk_in_reset.reset_n
	);

	wire          tristate_controller_tcm_chipselect_n_out;                                                                  // tristate_controller:tcm_chipselect_n_out -> tristate_conduit_pin_sharer:tcs0_chipselect_n_out
	wire          tristate_controller_tcm_grant;                                                                             // tristate_conduit_pin_sharer:tcs0_grant -> tristate_controller:tcm_grant
	wire          tristate_controller_tcm_data_outen;                                                                        // tristate_controller:tcm_data_outen -> tristate_conduit_pin_sharer:tcs0_data_outen
	wire          tristate_controller_tcm_byteenable_out;                                                                    // tristate_controller:tcm_byteenable_out -> tristate_conduit_pin_sharer:tcs0_byteenable_out
	wire          tristate_controller_tcm_request;                                                                           // tristate_controller:tcm_request -> tristate_conduit_pin_sharer:tcs0_request
	wire          tristate_controller_tcm_begintransfer_out;                                                                 // tristate_controller:tcm_begintransfer_out -> tristate_conduit_pin_sharer:tcs0_begintransfer_out
	wire    [7:0] tristate_controller_tcm_data_out;                                                                          // tristate_controller:tcm_data_out -> tristate_conduit_pin_sharer:tcs0_data_out
	wire          tristate_controller_tcm_write_n_out;                                                                       // tristate_controller:tcm_write_n_out -> tristate_conduit_pin_sharer:tcs0_write_n_out
	wire   [21:0] tristate_controller_tcm_address_out;                                                                       // tristate_controller:tcm_address_out -> tristate_conduit_pin_sharer:tcs0_address_out
	wire    [7:0] tristate_controller_tcm_data_in;                                                                           // tristate_conduit_pin_sharer:tcs0_data_in -> tristate_controller:tcm_data_in
	wire          tristate_controller_tcm_read_n_out;                                                                        // tristate_controller:tcm_read_n_out -> tristate_conduit_pin_sharer:tcs0_read_n_out
	wire    [0:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_byteenable_out_out;                                // tristate_conduit_pin_sharer:tristate_controller_tcm_byteenable_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_byteenable_out
	wire    [7:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_in;                                       // tristate_conduit_bridge:tcs_tristate_controller_tcm_data_in -> tristate_conduit_pin_sharer:tristate_controller_tcm_data_in
	wire    [0:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_read_n_out_out;                                    // tristate_conduit_pin_sharer:tristate_controller_tcm_read_n_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_read_n_out
	wire          tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_outen;                                    // tristate_conduit_pin_sharer:tristate_controller_tcm_data_outen -> tristate_conduit_bridge:tcs_tristate_controller_tcm_data_outen
	wire    [0:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_write_n_out_out;                                   // tristate_conduit_pin_sharer:tristate_controller_tcm_write_n_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_write_n_out
	wire          tristate_conduit_pin_sharer_tcm_grant;                                                                     // tristate_conduit_bridge:grant -> tristate_conduit_pin_sharer:grant
	wire    [0:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_begintransfer_out_out;                             // tristate_conduit_pin_sharer:tristate_controller_tcm_begintransfer_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_begintransfer_out
	wire          tristate_conduit_pin_sharer_tcm_request;                                                                   // tristate_conduit_pin_sharer:request -> tristate_conduit_bridge:request
	wire   [21:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_address_out_out;                                   // tristate_conduit_pin_sharer:tristate_controller_tcm_address_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_address_out
	wire    [7:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_out;                                      // tristate_conduit_pin_sharer:tristate_controller_tcm_data_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_data_out
	wire    [0:0] tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_chipselect_n_out_out;                              // tristate_conduit_pin_sharer:tristate_controller_tcm_chipselect_n_out -> tristate_conduit_bridge:tcs_tristate_controller_tcm_chipselect_n_out
	wire          main_pll_sys_clk_clk;                                                                                      // main_pll:sys_clk -> [add_button:clk, add_button_s1_translator:clk, add_button_s1_translator_avalon_universal_slave_0_agent:clk, add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, audio_config:clk, audio_config_avalon_av_config_slave_translator:clk, audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, barcode_scanner_ps2:clk, barcode_scanner_ps2_avalon_ps2_slave_translator:clk, barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:clk, barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, burst_adapter_004:clk, burst_adapter_005:clk, burst_adapter_006:clk, burst_adapter_007:clk, burst_adapter_008:clk, burst_adapter_009:clk, burst_adapter_010:clk, burst_adapter_011:clk, burst_adapter_012:clk, burst_adapter_013:clk, burst_adapter_014:clk, burst_adapter_016:clk, burst_adapter_017:clk, burst_adapter_018:clk, cancel_button:clk, cancel_button_s1_translator:clk, cancel_button_s1_translator_avalon_universal_slave_0_agent:clk, cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, character_lcd:clk, character_lcd_avalon_lcd_slave_translator:clk, character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_006:clk, cmd_xbar_mux_018:clk, crosser:in_clk, crosser_001:out_clk, dm9000a_if_ethernet:avs_s1_clk_iCLK, dm9000a_if_ethernet_s1_translator:clk, dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:clk, dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, green_leds:clk, green_leds_s1_translator:clk, green_leds_s1_translator_avalon_universal_slave_0_agent:clk, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, nios2_qsys:clk, nios2_qsys_data_master_translator:clk, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_instruction_master_translator:clk, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_jtag_debug_module_translator:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2:clk, onchip_memory2_s1_translator:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, red_leds:clk, red_leds_s1_translator:clk, red_leds_s1_translator_avalon_universal_slave_0_agent:clk, red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, remove_button:clk, remove_button_s1_translator:clk, remove_button_s1_translator_avalon_universal_slave_0_agent:clk, remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram:clk, sram_avalon_sram_slave_translator:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch:clk, switch_s1_translator:clk, switch_s1_translator_avalon_universal_slave_0_agent:clk, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys:clock, sysid_qsys_control_slave_translator:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, tristate_conduit_bridge:clk, tristate_conduit_pin_sharer:clk_clk, tristate_controller:clk_clk, tristate_controller_uas_translator:clk, tristate_controller_uas_translator_avalon_universal_slave_0_agent:clk, tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk]
	wire          main_pll_audio_clk_clk;                                                                                    // main_pll:AUD_CLK -> [audio_core:clk, audio_core_avalon_audio_slave_translator:clk, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:clk, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter_015:clk, crosser:out_clk, crosser_001:in_clk, id_router_015:clk, irq_synchronizer:receiver_clk, rsp_xbar_demux_015:clk, rst_controller_001:clk]
	wire    [3:0] nios2_qsys_data_master_burstcount;                                                                         // nios2_qsys:d_burstcount -> nios2_qsys_data_master_translator:av_burstcount
	wire          nios2_qsys_data_master_waitrequest;                                                                        // nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	wire   [31:0] nios2_qsys_data_master_writedata;                                                                          // nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	wire   [24:0] nios2_qsys_data_master_address;                                                                            // nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	wire          nios2_qsys_data_master_write;                                                                              // nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	wire          nios2_qsys_data_master_read;                                                                               // nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	wire   [31:0] nios2_qsys_data_master_readdata;                                                                           // nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	wire          nios2_qsys_data_master_debugaccess;                                                                        // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	wire          nios2_qsys_data_master_readdatavalid;                                                                      // nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	wire    [3:0] nios2_qsys_data_master_byteenable;                                                                         // nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	wire    [3:0] nios2_qsys_instruction_master_burstcount;                                                                  // nios2_qsys:i_burstcount -> nios2_qsys_instruction_master_translator:av_burstcount
	wire          nios2_qsys_instruction_master_waitrequest;                                                                 // nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	wire   [24:0] nios2_qsys_instruction_master_address;                                                                     // nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	wire          nios2_qsys_instruction_master_read;                                                                        // nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_instruction_master_readdata;                                                                    // nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	wire          nios2_qsys_instruction_master_readdatavalid;                                                               // nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                     // nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address;                                       // nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                    // nios2_qsys_jtag_debug_module_translator:av_chipselect -> nios2_qsys:jtag_debug_module_select
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write;                                         // nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                      // nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                 // nios2_qsys_jtag_debug_module_translator:av_begintransfer -> nios2_qsys:jtag_debug_module_begintransfer
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                   // nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                    // nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire          character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                 // character_lcd:waitrequest -> character_lcd_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                   // character_lcd_avalon_lcd_slave_translator:av_writedata -> character_lcd:writedata
	wire    [0:0] character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                     // character_lcd_avalon_lcd_slave_translator:av_address -> character_lcd:address
	wire          character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                  // character_lcd_avalon_lcd_slave_translator:av_chipselect -> character_lcd:chipselect
	wire          character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                       // character_lcd_avalon_lcd_slave_translator:av_write -> character_lcd:write
	wire          character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                        // character_lcd_avalon_lcd_slave_translator:av_read -> character_lcd:read
	wire    [7:0] character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                    // character_lcd:readdata -> character_lcd_avalon_lcd_slave_translator:av_readdata
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                           // sram_avalon_sram_slave_translator:av_writedata -> sram:writedata
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                             // sram_avalon_sram_slave_translator:av_address -> sram:address
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                               // sram_avalon_sram_slave_translator:av_write -> sram:write
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                // sram_avalon_sram_slave_translator:av_read -> sram:read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                            // sram:readdata -> sram_avalon_sram_slave_translator:av_readdata
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                       // sram:readdatavalid -> sram_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                          // sram_avalon_sram_slave_translator:av_byteenable -> sram:byteenable
	wire    [0:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_address;                                           // sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata;                                          // sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_writedata;                                                    // green_leds_s1_translator:av_writedata -> green_leds:writedata
	wire    [1:0] green_leds_s1_translator_avalon_anti_slave_0_address;                                                      // green_leds_s1_translator:av_address -> green_leds:address
	wire          green_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                   // green_leds_s1_translator:av_chipselect -> green_leds:chipselect
	wire          green_leds_s1_translator_avalon_anti_slave_0_write;                                                        // green_leds_s1_translator:av_write -> green_leds:write_n
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_readdata;                                                     // green_leds:readdata -> green_leds_s1_translator:av_readdata
	wire   [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_writedata;                                                // onchip_memory2_s1_translator:av_writedata -> onchip_memory2:writedata
	wire   [11:0] onchip_memory2_s1_translator_avalon_anti_slave_0_address;                                                  // onchip_memory2_s1_translator:av_address -> onchip_memory2:address
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect;                                               // onchip_memory2_s1_translator:av_chipselect -> onchip_memory2:chipselect
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_clken;                                                    // onchip_memory2_s1_translator:av_clken -> onchip_memory2:clken
	wire          onchip_memory2_s1_translator_avalon_anti_slave_0_write;                                                    // onchip_memory2_s1_translator:av_write -> onchip_memory2:write
	wire   [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_readdata;                                                 // onchip_memory2:readdata -> onchip_memory2_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable;                                               // onchip_memory2_s1_translator:av_byteenable -> onchip_memory2:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                       // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                         // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                           // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                        // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                             // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                              // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                          // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                     // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                        // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] switch_s1_translator_avalon_anti_slave_0_writedata;                                                        // switch_s1_translator:av_writedata -> switch:writedata
	wire    [1:0] switch_s1_translator_avalon_anti_slave_0_address;                                                          // switch_s1_translator:av_address -> switch:address
	wire          switch_s1_translator_avalon_anti_slave_0_chipselect;                                                       // switch_s1_translator:av_chipselect -> switch:chipselect
	wire          switch_s1_translator_avalon_anti_slave_0_write;                                                            // switch_s1_translator:av_write -> switch:write_n
	wire   [31:0] switch_s1_translator_avalon_anti_slave_0_readdata;                                                         // switch:readdata -> switch_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                         // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                           // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                                        // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                             // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                          // timer:readdata -> timer_s1_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                    // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                      // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                        // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                     // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                          // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                           // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                       // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] add_button_s1_translator_avalon_anti_slave_0_writedata;                                                    // add_button_s1_translator:av_writedata -> add_button:writedata
	wire    [1:0] add_button_s1_translator_avalon_anti_slave_0_address;                                                      // add_button_s1_translator:av_address -> add_button:address
	wire          add_button_s1_translator_avalon_anti_slave_0_chipselect;                                                   // add_button_s1_translator:av_chipselect -> add_button:chipselect
	wire          add_button_s1_translator_avalon_anti_slave_0_write;                                                        // add_button_s1_translator:av_write -> add_button:write_n
	wire   [31:0] add_button_s1_translator_avalon_anti_slave_0_readdata;                                                     // add_button:readdata -> add_button_s1_translator:av_readdata
	wire   [31:0] remove_button_s1_translator_avalon_anti_slave_0_writedata;                                                 // remove_button_s1_translator:av_writedata -> remove_button:writedata
	wire    [1:0] remove_button_s1_translator_avalon_anti_slave_0_address;                                                   // remove_button_s1_translator:av_address -> remove_button:address
	wire          remove_button_s1_translator_avalon_anti_slave_0_chipselect;                                                // remove_button_s1_translator:av_chipselect -> remove_button:chipselect
	wire          remove_button_s1_translator_avalon_anti_slave_0_write;                                                     // remove_button_s1_translator:av_write -> remove_button:write_n
	wire   [31:0] remove_button_s1_translator_avalon_anti_slave_0_readdata;                                                  // remove_button:readdata -> remove_button_s1_translator:av_readdata
	wire   [31:0] cancel_button_s1_translator_avalon_anti_slave_0_writedata;                                                 // cancel_button_s1_translator:av_writedata -> cancel_button:writedata
	wire    [1:0] cancel_button_s1_translator_avalon_anti_slave_0_address;                                                   // cancel_button_s1_translator:av_address -> cancel_button:address
	wire          cancel_button_s1_translator_avalon_anti_slave_0_chipselect;                                                // cancel_button_s1_translator:av_chipselect -> cancel_button:chipselect
	wire          cancel_button_s1_translator_avalon_anti_slave_0_write;                                                     // cancel_button_s1_translator:av_write -> cancel_button:write_n
	wire   [31:0] cancel_button_s1_translator_avalon_anti_slave_0_readdata;                                                  // cancel_button:readdata -> cancel_button_s1_translator:av_readdata
	wire   [31:0] red_leds_s1_translator_avalon_anti_slave_0_writedata;                                                      // red_leds_s1_translator:av_writedata -> red_leds:writedata
	wire    [1:0] red_leds_s1_translator_avalon_anti_slave_0_address;                                                        // red_leds_s1_translator:av_address -> red_leds:address
	wire          red_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                     // red_leds_s1_translator:av_chipselect -> red_leds:chipselect
	wire          red_leds_s1_translator_avalon_anti_slave_0_write;                                                          // red_leds_s1_translator:av_write -> red_leds:write_n
	wire   [31:0] red_leds_s1_translator_avalon_anti_slave_0_readdata;                                                       // red_leds:readdata -> red_leds_s1_translator:av_readdata
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest;                           // barcode_scanner_ps2:waitrequest -> barcode_scanner_ps2_avalon_ps2_slave_translator:av_waitrequest
	wire   [31:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata;                             // barcode_scanner_ps2_avalon_ps2_slave_translator:av_writedata -> barcode_scanner_ps2:writedata
	wire    [0:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_address;                               // barcode_scanner_ps2_avalon_ps2_slave_translator:av_address -> barcode_scanner_ps2:address
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect;                            // barcode_scanner_ps2_avalon_ps2_slave_translator:av_chipselect -> barcode_scanner_ps2:chipselect
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_write;                                 // barcode_scanner_ps2_avalon_ps2_slave_translator:av_write -> barcode_scanner_ps2:write
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_read;                                  // barcode_scanner_ps2_avalon_ps2_slave_translator:av_read -> barcode_scanner_ps2:read
	wire   [31:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata;                              // barcode_scanner_ps2:readdata -> barcode_scanner_ps2_avalon_ps2_slave_translator:av_readdata
	wire    [3:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable;                            // barcode_scanner_ps2_avalon_ps2_slave_translator:av_byteenable -> barcode_scanner_ps2:byteenable
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_writedata;                                    // audio_core_avalon_audio_slave_translator:av_writedata -> audio_core:writedata
	wire    [1:0] audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_address;                                      // audio_core_avalon_audio_slave_translator:av_address -> audio_core:address
	wire          audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect;                                   // audio_core_avalon_audio_slave_translator:av_chipselect -> audio_core:chipselect
	wire          audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_write;                                        // audio_core_avalon_audio_slave_translator:av_write -> audio_core:write
	wire          audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_read;                                         // audio_core_avalon_audio_slave_translator:av_read -> audio_core:read
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_readdata;                                     // audio_core:readdata -> audio_core_avalon_audio_slave_translator:av_readdata
	wire          audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                            // audio_config:waitrequest -> audio_config_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                              // audio_config_avalon_av_config_slave_translator:av_writedata -> audio_config:writedata
	wire    [1:0] audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                                // audio_config_avalon_av_config_slave_translator:av_address -> audio_config:address
	wire          audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                  // audio_config_avalon_av_config_slave_translator:av_write -> audio_config:write
	wire          audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                   // audio_config_avalon_av_config_slave_translator:av_read -> audio_config:read
	wire   [31:0] audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                               // audio_config:readdata -> audio_config_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                             // audio_config_avalon_av_config_slave_translator:av_byteenable -> audio_config:byteenable
	wire   [15:0] dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_writedata;                                           // dm9000a_if_ethernet_s1_translator:av_writedata -> dm9000a_if_ethernet:avs_s1_writedata_iDATA
	wire    [0:0] dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_address;                                             // dm9000a_if_ethernet_s1_translator:av_address -> dm9000a_if_ethernet:avs_s1_address_iCMD
	wire          dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_chipselect;                                          // dm9000a_if_ethernet_s1_translator:av_chipselect -> dm9000a_if_ethernet:avs_s1_chipselect_n_iCS_N
	wire          dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_write;                                               // dm9000a_if_ethernet_s1_translator:av_write -> dm9000a_if_ethernet:avs_s1_write_n_iWR_N
	wire          dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_read;                                                // dm9000a_if_ethernet_s1_translator:av_read -> dm9000a_if_ethernet:avs_s1_read_n_iRD_N
	wire   [15:0] dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_readdata;                                            // dm9000a_if_ethernet:avs_s1_readdata_oDATA -> dm9000a_if_ethernet_s1_translator:av_readdata
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_waitrequest;                                        // tristate_controller:uas_waitrequest -> tristate_controller_uas_translator:av_waitrequest
	wire    [0:0] tristate_controller_uas_translator_avalon_anti_slave_0_burstcount;                                         // tristate_controller_uas_translator:av_burstcount -> tristate_controller:uas_burstcount
	wire    [7:0] tristate_controller_uas_translator_avalon_anti_slave_0_writedata;                                          // tristate_controller_uas_translator:av_writedata -> tristate_controller:uas_writedata
	wire   [21:0] tristate_controller_uas_translator_avalon_anti_slave_0_address;                                            // tristate_controller_uas_translator:av_address -> tristate_controller:uas_address
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_lock;                                               // tristate_controller_uas_translator:av_lock -> tristate_controller:uas_lock
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_write;                                              // tristate_controller_uas_translator:av_write -> tristate_controller:uas_write
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_read;                                               // tristate_controller_uas_translator:av_read -> tristate_controller:uas_read
	wire    [7:0] tristate_controller_uas_translator_avalon_anti_slave_0_readdata;                                           // tristate_controller:uas_readdata -> tristate_controller_uas_translator:av_readdata
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_debugaccess;                                        // tristate_controller_uas_translator:av_debugaccess -> tristate_controller:uas_debugaccess
	wire          tristate_controller_uas_translator_avalon_anti_slave_0_readdatavalid;                                      // tristate_controller:uas_readdatavalid -> tristate_controller_uas_translator:av_readdatavalid
	wire    [0:0] tristate_controller_uas_translator_avalon_anti_slave_0_byteenable;                                         // tristate_controller_uas_translator:av_byteenable -> tristate_controller:uas_byteenable
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest;                                   // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	wire    [5:0] nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount;                                    // nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_writedata;                                     // nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] nios2_qsys_data_master_translator_avalon_universal_master_0_address;                                       // nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_lock;                                          // nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_write;                                         // nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_read;                                          // nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_readdata;                                      // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess;                                   // nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable;                                    // nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid;                                 // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest;                            // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	wire    [5:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount;                             // nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata;                              // nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_address;                                // nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock;                                   // nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_write;                                  // nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_read;                                   // nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata;                               // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess;                            // nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable;                             // nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid;                          // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	wire   [24:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                        // nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // character_lcd_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_avalon_lcd_slave_translator:uav_writedata
	wire   [24:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // character_lcd_avalon_lcd_slave_translator:uav_readdata -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // character_lcd_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_avalon_lcd_slave_translator:uav_debugaccess
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // sram_avalon_sram_slave_translator:uav_waitrequest -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_avalon_sram_slave_translator:uav_writedata
	wire   [24:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_avalon_sram_slave_translator:uav_address
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_avalon_sram_slave_translator:uav_write
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_avalon_sram_slave_translator:uav_lock
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // sram_avalon_sram_slave_translator:uav_readdata -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // sram_avalon_sram_slave_translator:uav_readdatavalid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_avalon_sram_slave_translator:uav_byteenable
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [90:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [90:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	wire   [24:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // green_leds_s1_translator:uav_waitrequest -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_leds_s1_translator:uav_burstcount
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_leds_s1_translator:uav_writedata
	wire   [24:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_leds_s1_translator:uav_address
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_leds_s1_translator:uav_write
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_leds_s1_translator:uav_lock
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_leds_s1_translator:uav_read
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // green_leds_s1_translator:uav_readdata -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // green_leds_s1_translator:uav_readdatavalid -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_leds_s1_translator:uav_debugaccess
	wire    [3:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_leds_s1_translator:uav_byteenable
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // onchip_memory2_s1_translator:uav_waitrequest -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_s1_translator:uav_writedata
	wire   [24:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_s1_translator:uav_address
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_s1_translator:uav_write
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_s1_translator:uav_lock
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_s1_translator:uav_read
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // onchip_memory2_s1_translator:uav_readdata -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // onchip_memory2_s1_translator:uav_readdatavalid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_s1_translator:uav_byteenable
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [24:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [90:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [90:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // switch_s1_translator:uav_waitrequest -> switch_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_s1_translator:uav_burstcount
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // switch_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_s1_translator:uav_writedata
	wire   [24:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // switch_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_s1_translator:uav_address
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // switch_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_s1_translator:uav_write
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // switch_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_s1_translator:uav_lock
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // switch_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_s1_translator:uav_read
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // switch_s1_translator:uav_readdata -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // switch_s1_translator:uav_readdatavalid -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // switch_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_s1_translator:uav_debugaccess
	wire    [3:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_s1_translator:uav_byteenable
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire   [24:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [24:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // add_button_s1_translator:uav_waitrequest -> add_button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] add_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // add_button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> add_button_s1_translator:uav_burstcount
	wire   [31:0] add_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // add_button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> add_button_s1_translator:uav_writedata
	wire   [24:0] add_button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // add_button_s1_translator_avalon_universal_slave_0_agent:m0_address -> add_button_s1_translator:uav_address
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // add_button_s1_translator_avalon_universal_slave_0_agent:m0_write -> add_button_s1_translator:uav_write
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // add_button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> add_button_s1_translator:uav_lock
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // add_button_s1_translator_avalon_universal_slave_0_agent:m0_read -> add_button_s1_translator:uav_read
	wire   [31:0] add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // add_button_s1_translator:uav_readdata -> add_button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // add_button_s1_translator:uav_readdatavalid -> add_button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // add_button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> add_button_s1_translator:uav_debugaccess
	wire    [3:0] add_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // add_button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> add_button_s1_translator:uav_byteenable
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // add_button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // add_button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // add_button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // add_button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> add_button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> add_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> add_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // add_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> add_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // remove_button_s1_translator:uav_waitrequest -> remove_button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] remove_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> remove_button_s1_translator:uav_burstcount
	wire   [31:0] remove_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> remove_button_s1_translator:uav_writedata
	wire   [24:0] remove_button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_address -> remove_button_s1_translator:uav_address
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_write -> remove_button_s1_translator:uav_write
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> remove_button_s1_translator:uav_lock
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_read -> remove_button_s1_translator:uav_read
	wire   [31:0] remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // remove_button_s1_translator:uav_readdata -> remove_button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // remove_button_s1_translator:uav_readdatavalid -> remove_button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> remove_button_s1_translator:uav_debugaccess
	wire    [3:0] remove_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // remove_button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> remove_button_s1_translator:uav_byteenable
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // remove_button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // remove_button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // remove_button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // remove_button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> remove_button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> remove_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> remove_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // remove_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> remove_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // cancel_button_s1_translator:uav_waitrequest -> cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> cancel_button_s1_translator:uav_burstcount
	wire   [31:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> cancel_button_s1_translator:uav_writedata
	wire   [24:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_address -> cancel_button_s1_translator:uav_address
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_write -> cancel_button_s1_translator:uav_write
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> cancel_button_s1_translator:uav_lock
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_read -> cancel_button_s1_translator:uav_read
	wire   [31:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // cancel_button_s1_translator:uav_readdata -> cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // cancel_button_s1_translator:uav_readdatavalid -> cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cancel_button_s1_translator:uav_debugaccess
	wire    [3:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // cancel_button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> cancel_button_s1_translator:uav_byteenable
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // cancel_button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // red_leds_s1_translator:uav_waitrequest -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> red_leds_s1_translator:uav_burstcount
	wire   [31:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> red_leds_s1_translator:uav_writedata
	wire   [24:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> red_leds_s1_translator:uav_address
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> red_leds_s1_translator:uav_write
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> red_leds_s1_translator:uav_lock
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> red_leds_s1_translator:uav_read
	wire   [31:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // red_leds_s1_translator:uav_readdata -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // red_leds_s1_translator:uav_readdatavalid -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> red_leds_s1_translator:uav_debugaccess
	wire    [3:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> red_leds_s1_translator:uav_byteenable
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // barcode_scanner_ps2_avalon_ps2_slave_translator:uav_waitrequest -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_burstcount
	wire   [31:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_writedata
	wire   [24:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_address -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_address
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_write -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_write
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_lock -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_lock
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_read -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_read
	wire   [31:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // barcode_scanner_ps2_avalon_ps2_slave_translator:uav_readdata -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // barcode_scanner_ps2_avalon_ps2_slave_translator:uav_readdatavalid -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_debugaccess
	wire    [3:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> barcode_scanner_ps2_avalon_ps2_slave_translator:uav_byteenable
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // audio_core_avalon_audio_slave_translator:uav_waitrequest -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_core_avalon_audio_slave_translator:uav_burstcount
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_core_avalon_audio_slave_translator:uav_writedata
	wire   [24:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_core_avalon_audio_slave_translator:uav_address
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_core_avalon_audio_slave_translator:uav_write
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_core_avalon_audio_slave_translator:uav_lock
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_core_avalon_audio_slave_translator:uav_read
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // audio_core_avalon_audio_slave_translator:uav_readdata -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // audio_core_avalon_audio_slave_translator:uav_readdatavalid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_core_avalon_audio_slave_translator:uav_debugaccess
	wire    [3:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_core_avalon_audio_slave_translator:uav_byteenable
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // audio_config_avalon_av_config_slave_translator:uav_waitrequest -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_config_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_config_avalon_av_config_slave_translator:uav_writedata
	wire   [24:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_config_avalon_av_config_slave_translator:uav_address
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_config_avalon_av_config_slave_translator:uav_write
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_config_avalon_av_config_slave_translator:uav_lock
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_config_avalon_av_config_slave_translator:uav_read
	wire   [31:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // audio_config_avalon_av_config_slave_translator:uav_readdata -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // audio_config_avalon_av_config_slave_translator:uav_readdatavalid -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_config_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_config_avalon_av_config_slave_translator:uav_byteenable
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // dm9000a_if_ethernet_s1_translator:uav_waitrequest -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dm9000a_if_ethernet_s1_translator:uav_burstcount
	wire   [31:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dm9000a_if_ethernet_s1_translator:uav_writedata
	wire   [24:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_address -> dm9000a_if_ethernet_s1_translator:uav_address
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_write -> dm9000a_if_ethernet_s1_translator:uav_write
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dm9000a_if_ethernet_s1_translator:uav_lock
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_read -> dm9000a_if_ethernet_s1_translator:uav_read
	wire   [31:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // dm9000a_if_ethernet_s1_translator:uav_readdata -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // dm9000a_if_ethernet_s1_translator:uav_readdatavalid -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dm9000a_if_ethernet_s1_translator:uav_debugaccess
	wire    [3:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dm9000a_if_ethernet_s1_translator:uav_byteenable
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // tristate_controller_uas_translator:uav_waitrequest -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> tristate_controller_uas_translator:uav_burstcount
	wire    [7:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                            // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> tristate_controller_uas_translator:uav_writedata
	wire   [24:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_address;                              // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_address -> tristate_controller_uas_translator:uav_address
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_write;                                // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_write -> tristate_controller_uas_translator:uav_write
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                 // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_lock -> tristate_controller_uas_translator:uav_lock
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_read;                                 // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_read -> tristate_controller_uas_translator:uav_read
	wire    [7:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                             // tristate_controller_uas_translator:uav_readdata -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // tristate_controller_uas_translator:uav_readdatavalid -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tristate_controller_uas_translator:uav_debugaccess
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // tristate_controller_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> tristate_controller_uas_translator:uav_byteenable
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                          // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [107:0] nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data;                                 // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                         // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [107:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                          // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_001:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [107:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [80:0] character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_001:sink_ready -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [89:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_002:sink_ready -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [107:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_003:sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [107:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_004:sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [107:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_005:sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_006:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // switch_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // switch_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // switch_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [107:0] switch_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // switch_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_007:sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [107:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_008:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_009:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // add_button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // add_button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // add_button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [107:0] add_button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // add_button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          add_button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_010:sink_ready -> add_button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // remove_button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // remove_button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // remove_button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [107:0] remove_button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // remove_button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          remove_button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_011:sink_ready -> remove_button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // cancel_button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // cancel_button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // cancel_button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [107:0] cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // cancel_button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> cancel_button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [107:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_013:sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [107:0] barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_014:sink_ready -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [107:0] audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_015:sink_ready -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [107:0] audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_016:sink_ready -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [107:0] dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_017:sink_ready -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [80:0] tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_data;                                 // tristate_controller_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_018:sink_ready -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                               // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                     // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                             // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [107:0] addr_router_src_data;                                                                                      // addr_router:src_data -> limiter:cmd_sink_data
	wire   [18:0] addr_router_src_channel;                                                                                   // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                     // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                               // limiter:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                     // limiter:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                             // limiter:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] limiter_rsp_src_data;                                                                                      // limiter:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_rsp_src_channel;                                                                                   // limiter:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                     // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                           // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                 // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                         // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [107:0] addr_router_001_src_data;                                                                                  // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [18:0] addr_router_001_src_channel;                                                                               // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                 // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                           // limiter_001:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                 // limiter_001:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                         // limiter_001:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] limiter_001_rsp_src_data;                                                                                  // limiter_001:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_001_rsp_src_channel;                                                                               // limiter_001:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                 // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                         // burst_adapter:source0_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                               // burst_adapter:source0_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                       // burst_adapter:source0_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_source0_data;                                                                                // burst_adapter:source0_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [18:0] burst_adapter_source0_channel;                                                                             // burst_adapter:source0_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                     // burst_adapter_001:source0_endofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                           // burst_adapter_001:source0_valid -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                   // burst_adapter_001:source0_startofpacket -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] burst_adapter_001_source0_data;                                                                            // burst_adapter_001:source0_data -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                           // character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [18:0] burst_adapter_001_source0_channel;                                                                         // burst_adapter_001:source0_channel -> character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                     // burst_adapter_002:source0_endofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                           // burst_adapter_002:source0_valid -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                   // burst_adapter_002:source0_startofpacket -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [89:0] burst_adapter_002_source0_data;                                                                            // burst_adapter_002:source0_data -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                           // sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [18:0] burst_adapter_002_source0_channel;                                                                         // burst_adapter_002:source0_channel -> sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                     // burst_adapter_003:source0_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                           // burst_adapter_003:source0_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                   // burst_adapter_003:source0_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_003_source0_data;                                                                            // burst_adapter_003:source0_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [18:0] burst_adapter_003_source0_channel;                                                                         // burst_adapter_003:source0_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                                     // burst_adapter_004:source0_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                           // burst_adapter_004:source0_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                                   // burst_adapter_004:source0_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_004_source0_data;                                                                            // burst_adapter_004:source0_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire   [18:0] burst_adapter_004_source0_channel;                                                                         // burst_adapter_004:source0_channel -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_005_source0_endofpacket;                                                                     // burst_adapter_005:source0_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_005_source0_valid;                                                                           // burst_adapter_005:source0_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_005_source0_startofpacket;                                                                   // burst_adapter_005:source0_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_005_source0_data;                                                                            // burst_adapter_005:source0_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_005_source0_ready;                                                                           // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_005:source0_ready
	wire   [18:0] burst_adapter_005_source0_channel;                                                                         // burst_adapter_005:source0_channel -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_006_source0_endofpacket;                                                                     // burst_adapter_006:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_006_source0_valid;                                                                           // burst_adapter_006:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_006_source0_startofpacket;                                                                   // burst_adapter_006:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [89:0] burst_adapter_006_source0_data;                                                                            // burst_adapter_006:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_006_source0_ready;                                                                           // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_006:source0_ready
	wire   [18:0] burst_adapter_006_source0_channel;                                                                         // burst_adapter_006:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_007_source0_endofpacket;                                                                     // burst_adapter_007:source0_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_007_source0_valid;                                                                           // burst_adapter_007:source0_valid -> switch_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_007_source0_startofpacket;                                                                   // burst_adapter_007:source0_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_007_source0_data;                                                                            // burst_adapter_007:source0_data -> switch_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_007_source0_ready;                                                                           // switch_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_007:source0_ready
	wire   [18:0] burst_adapter_007_source0_channel;                                                                         // burst_adapter_007:source0_channel -> switch_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_008_source0_endofpacket;                                                                     // burst_adapter_008:source0_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_008_source0_valid;                                                                           // burst_adapter_008:source0_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_008_source0_startofpacket;                                                                   // burst_adapter_008:source0_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_008_source0_data;                                                                            // burst_adapter_008:source0_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_008_source0_ready;                                                                           // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_008:source0_ready
	wire   [18:0] burst_adapter_008_source0_channel;                                                                         // burst_adapter_008:source0_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_009_source0_endofpacket;                                                                     // burst_adapter_009:source0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_009_source0_valid;                                                                           // burst_adapter_009:source0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_009_source0_startofpacket;                                                                   // burst_adapter_009:source0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_009_source0_data;                                                                            // burst_adapter_009:source0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_009_source0_ready;                                                                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_009:source0_ready
	wire   [18:0] burst_adapter_009_source0_channel;                                                                         // burst_adapter_009:source0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_010_source0_endofpacket;                                                                     // burst_adapter_010:source0_endofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_010_source0_valid;                                                                           // burst_adapter_010:source0_valid -> add_button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_010_source0_startofpacket;                                                                   // burst_adapter_010:source0_startofpacket -> add_button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_010_source0_data;                                                                            // burst_adapter_010:source0_data -> add_button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_010_source0_ready;                                                                           // add_button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_010:source0_ready
	wire   [18:0] burst_adapter_010_source0_channel;                                                                         // burst_adapter_010:source0_channel -> add_button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_011_source0_endofpacket;                                                                     // burst_adapter_011:source0_endofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_011_source0_valid;                                                                           // burst_adapter_011:source0_valid -> remove_button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_011_source0_startofpacket;                                                                   // burst_adapter_011:source0_startofpacket -> remove_button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_011_source0_data;                                                                            // burst_adapter_011:source0_data -> remove_button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_011_source0_ready;                                                                           // remove_button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_011:source0_ready
	wire   [18:0] burst_adapter_011_source0_channel;                                                                         // burst_adapter_011:source0_channel -> remove_button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_012_source0_endofpacket;                                                                     // burst_adapter_012:source0_endofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_012_source0_valid;                                                                           // burst_adapter_012:source0_valid -> cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_012_source0_startofpacket;                                                                   // burst_adapter_012:source0_startofpacket -> cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_012_source0_data;                                                                            // burst_adapter_012:source0_data -> cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_012_source0_ready;                                                                           // cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_012:source0_ready
	wire   [18:0] burst_adapter_012_source0_channel;                                                                         // burst_adapter_012:source0_channel -> cancel_button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_013_source0_endofpacket;                                                                     // burst_adapter_013:source0_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_013_source0_valid;                                                                           // burst_adapter_013:source0_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_013_source0_startofpacket;                                                                   // burst_adapter_013:source0_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_013_source0_data;                                                                            // burst_adapter_013:source0_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_013_source0_ready;                                                                           // red_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_013:source0_ready
	wire   [18:0] burst_adapter_013_source0_channel;                                                                         // burst_adapter_013:source0_channel -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_014_source0_endofpacket;                                                                     // burst_adapter_014:source0_endofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_014_source0_valid;                                                                           // burst_adapter_014:source0_valid -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_014_source0_startofpacket;                                                                   // burst_adapter_014:source0_startofpacket -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_014_source0_data;                                                                            // burst_adapter_014:source0_data -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_014_source0_ready;                                                                           // barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_014:source0_ready
	wire   [18:0] burst_adapter_014_source0_channel;                                                                         // burst_adapter_014:source0_channel -> barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_015_source0_endofpacket;                                                                     // burst_adapter_015:source0_endofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_015_source0_valid;                                                                           // burst_adapter_015:source0_valid -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_015_source0_startofpacket;                                                                   // burst_adapter_015:source0_startofpacket -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_015_source0_data;                                                                            // burst_adapter_015:source0_data -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_015_source0_ready;                                                                           // audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_015:source0_ready
	wire   [18:0] burst_adapter_015_source0_channel;                                                                         // burst_adapter_015:source0_channel -> audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_016_source0_endofpacket;                                                                     // burst_adapter_016:source0_endofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_016_source0_valid;                                                                           // burst_adapter_016:source0_valid -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_016_source0_startofpacket;                                                                   // burst_adapter_016:source0_startofpacket -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_016_source0_data;                                                                            // burst_adapter_016:source0_data -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_016_source0_ready;                                                                           // audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_016:source0_ready
	wire   [18:0] burst_adapter_016_source0_channel;                                                                         // burst_adapter_016:source0_channel -> audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_017_source0_endofpacket;                                                                     // burst_adapter_017:source0_endofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_017_source0_valid;                                                                           // burst_adapter_017:source0_valid -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_017_source0_startofpacket;                                                                   // burst_adapter_017:source0_startofpacket -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_017_source0_data;                                                                            // burst_adapter_017:source0_data -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_017_source0_ready;                                                                           // dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_017:source0_ready
	wire   [18:0] burst_adapter_017_source0_channel;                                                                         // burst_adapter_017:source0_channel -> dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_018_source0_endofpacket;                                                                     // burst_adapter_018:source0_endofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_018_source0_valid;                                                                           // burst_adapter_018:source0_valid -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_018_source0_startofpacket;                                                                   // burst_adapter_018:source0_startofpacket -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] burst_adapter_018_source0_data;                                                                            // burst_adapter_018:source0_data -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_018_source0_ready;                                                                           // tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_018:source0_ready
	wire   [18:0] burst_adapter_018_source0_channel;                                                                         // burst_adapter_018:source0_channel -> tristate_controller_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                            // rst_controller:reset_out -> [add_button:reset_n, add_button_s1_translator:reset, add_button_s1_translator_avalon_universal_slave_0_agent:reset, add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, audio_config:reset, audio_config_avalon_av_config_slave_translator:reset, audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, barcode_scanner_ps2:reset, barcode_scanner_ps2_avalon_ps2_slave_translator:reset, barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:reset, barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, burst_adapter_004:reset, burst_adapter_005:reset, burst_adapter_006:reset, burst_adapter_007:reset, burst_adapter_008:reset, burst_adapter_009:reset, burst_adapter_010:reset, burst_adapter_011:reset, burst_adapter_012:reset, burst_adapter_013:reset, burst_adapter_014:reset, burst_adapter_016:reset, burst_adapter_017:reset, burst_adapter_018:reset, cancel_button:reset_n, cancel_button_s1_translator:reset, cancel_button_s1_translator_avalon_universal_slave_0_agent:reset, cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, character_lcd:reset, character_lcd_avalon_lcd_slave_translator:reset, character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_018:reset, crosser:in_reset, crosser_001:out_reset, dm9000a_if_ethernet:avs_s1_reset_n_iRST_N, dm9000a_if_ethernet_s1_translator:reset, dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent:reset, dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, green_leds:reset_n, green_leds_s1_translator:reset, green_leds_s1_translator_avalon_universal_slave_0_agent:reset, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys:reset_n, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2:reset, onchip_memory2_s1_translator:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, red_leds:reset_n, red_leds_s1_translator:reset, red_leds_s1_translator_avalon_universal_slave_0_agent:reset, red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, remove_button:reset_n, remove_button_s1_translator:reset, remove_button_s1_translator_avalon_universal_slave_0_agent:reset, remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram:reset, sram_avalon_sram_slave_translator:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch:reset_n, switch_s1_translator:reset, switch_s1_translator_avalon_universal_slave_0_agent:reset, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys:reset_n, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tristate_conduit_bridge:reset, tristate_conduit_pin_sharer:reset_reset, tristate_controller:reset_reset, tristate_controller_uas_translator:reset, tristate_controller_uas_translator_avalon_universal_slave_0_agent:reset, tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire          nios2_qsys_jtag_debug_module_reset_reset;                                                                  // nios2_qsys:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire          main_pll_sys_clk_reset_reset;                                                                              // main_pll:sys_reset_n -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2]
	wire          rst_controller_001_reset_out_reset;                                                                        // rst_controller_001:reset_out -> [audio_core:reset, audio_core_avalon_audio_slave_translator:reset, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent:reset, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_015:reset, crosser:out_reset, crosser_001:in_reset, id_router_015:reset, irq_synchronizer:receiver_reset, rsp_xbar_demux_015:reset]
	wire          rst_controller_002_reset_out_reset;                                                                        // rst_controller_002:reset_out -> main_pll:reset
	wire          cmd_xbar_demux_src0_endofpacket;                                                                           // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                 // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                         // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src0_data;                                                                                  // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [18:0] cmd_xbar_demux_src0_channel;                                                                               // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                 // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                           // cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                 // cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                         // cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	wire  [107:0] cmd_xbar_demux_src1_data;                                                                                  // cmd_xbar_demux:src1_data -> width_adapter:in_data
	wire   [18:0] cmd_xbar_demux_src1_channel;                                                                               // cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                           // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                 // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                         // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src2_data;                                                                                  // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [18:0] cmd_xbar_demux_src2_channel;                                                                               // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                 // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                           // cmd_xbar_demux:src3_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                 // cmd_xbar_demux:src3_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                         // cmd_xbar_demux:src3_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src3_data;                                                                                  // cmd_xbar_demux:src3_data -> burst_adapter_003:sink0_data
	wire   [18:0] cmd_xbar_demux_src3_channel;                                                                               // cmd_xbar_demux:src3_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_demux_src4_endofpacket;                                                                           // cmd_xbar_demux:src4_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                 // cmd_xbar_demux:src4_valid -> burst_adapter_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                         // cmd_xbar_demux:src4_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src4_data;                                                                                  // cmd_xbar_demux:src4_data -> burst_adapter_004:sink0_data
	wire   [18:0] cmd_xbar_demux_src4_channel;                                                                               // cmd_xbar_demux:src4_channel -> burst_adapter_004:sink0_channel
	wire          cmd_xbar_demux_src5_endofpacket;                                                                           // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                 // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                         // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src5_data;                                                                                  // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [18:0] cmd_xbar_demux_src5_channel;                                                                               // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                 // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire          cmd_xbar_demux_src6_endofpacket;                                                                           // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                                 // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                         // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src6_data;                                                                                  // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [18:0] cmd_xbar_demux_src6_channel;                                                                               // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_src6_ready;                                                                                 // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire          cmd_xbar_demux_src7_endofpacket;                                                                           // cmd_xbar_demux:src7_endofpacket -> burst_adapter_007:sink0_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                                 // cmd_xbar_demux:src7_valid -> burst_adapter_007:sink0_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                         // cmd_xbar_demux:src7_startofpacket -> burst_adapter_007:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src7_data;                                                                                  // cmd_xbar_demux:src7_data -> burst_adapter_007:sink0_data
	wire   [18:0] cmd_xbar_demux_src7_channel;                                                                               // cmd_xbar_demux:src7_channel -> burst_adapter_007:sink0_channel
	wire          cmd_xbar_demux_src8_endofpacket;                                                                           // cmd_xbar_demux:src8_endofpacket -> burst_adapter_008:sink0_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                                 // cmd_xbar_demux:src8_valid -> burst_adapter_008:sink0_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                         // cmd_xbar_demux:src8_startofpacket -> burst_adapter_008:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src8_data;                                                                                  // cmd_xbar_demux:src8_data -> burst_adapter_008:sink0_data
	wire   [18:0] cmd_xbar_demux_src8_channel;                                                                               // cmd_xbar_demux:src8_channel -> burst_adapter_008:sink0_channel
	wire          cmd_xbar_demux_src9_endofpacket;                                                                           // cmd_xbar_demux:src9_endofpacket -> burst_adapter_009:sink0_endofpacket
	wire          cmd_xbar_demux_src9_valid;                                                                                 // cmd_xbar_demux:src9_valid -> burst_adapter_009:sink0_valid
	wire          cmd_xbar_demux_src9_startofpacket;                                                                         // cmd_xbar_demux:src9_startofpacket -> burst_adapter_009:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src9_data;                                                                                  // cmd_xbar_demux:src9_data -> burst_adapter_009:sink0_data
	wire   [18:0] cmd_xbar_demux_src9_channel;                                                                               // cmd_xbar_demux:src9_channel -> burst_adapter_009:sink0_channel
	wire          cmd_xbar_demux_src10_endofpacket;                                                                          // cmd_xbar_demux:src10_endofpacket -> burst_adapter_010:sink0_endofpacket
	wire          cmd_xbar_demux_src10_valid;                                                                                // cmd_xbar_demux:src10_valid -> burst_adapter_010:sink0_valid
	wire          cmd_xbar_demux_src10_startofpacket;                                                                        // cmd_xbar_demux:src10_startofpacket -> burst_adapter_010:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src10_data;                                                                                 // cmd_xbar_demux:src10_data -> burst_adapter_010:sink0_data
	wire   [18:0] cmd_xbar_demux_src10_channel;                                                                              // cmd_xbar_demux:src10_channel -> burst_adapter_010:sink0_channel
	wire          cmd_xbar_demux_src11_endofpacket;                                                                          // cmd_xbar_demux:src11_endofpacket -> burst_adapter_011:sink0_endofpacket
	wire          cmd_xbar_demux_src11_valid;                                                                                // cmd_xbar_demux:src11_valid -> burst_adapter_011:sink0_valid
	wire          cmd_xbar_demux_src11_startofpacket;                                                                        // cmd_xbar_demux:src11_startofpacket -> burst_adapter_011:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src11_data;                                                                                 // cmd_xbar_demux:src11_data -> burst_adapter_011:sink0_data
	wire   [18:0] cmd_xbar_demux_src11_channel;                                                                              // cmd_xbar_demux:src11_channel -> burst_adapter_011:sink0_channel
	wire          cmd_xbar_demux_src12_endofpacket;                                                                          // cmd_xbar_demux:src12_endofpacket -> burst_adapter_012:sink0_endofpacket
	wire          cmd_xbar_demux_src12_valid;                                                                                // cmd_xbar_demux:src12_valid -> burst_adapter_012:sink0_valid
	wire          cmd_xbar_demux_src12_startofpacket;                                                                        // cmd_xbar_demux:src12_startofpacket -> burst_adapter_012:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src12_data;                                                                                 // cmd_xbar_demux:src12_data -> burst_adapter_012:sink0_data
	wire   [18:0] cmd_xbar_demux_src12_channel;                                                                              // cmd_xbar_demux:src12_channel -> burst_adapter_012:sink0_channel
	wire          cmd_xbar_demux_src13_endofpacket;                                                                          // cmd_xbar_demux:src13_endofpacket -> burst_adapter_013:sink0_endofpacket
	wire          cmd_xbar_demux_src13_valid;                                                                                // cmd_xbar_demux:src13_valid -> burst_adapter_013:sink0_valid
	wire          cmd_xbar_demux_src13_startofpacket;                                                                        // cmd_xbar_demux:src13_startofpacket -> burst_adapter_013:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src13_data;                                                                                 // cmd_xbar_demux:src13_data -> burst_adapter_013:sink0_data
	wire   [18:0] cmd_xbar_demux_src13_channel;                                                                              // cmd_xbar_demux:src13_channel -> burst_adapter_013:sink0_channel
	wire          cmd_xbar_demux_src14_endofpacket;                                                                          // cmd_xbar_demux:src14_endofpacket -> burst_adapter_014:sink0_endofpacket
	wire          cmd_xbar_demux_src14_valid;                                                                                // cmd_xbar_demux:src14_valid -> burst_adapter_014:sink0_valid
	wire          cmd_xbar_demux_src14_startofpacket;                                                                        // cmd_xbar_demux:src14_startofpacket -> burst_adapter_014:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src14_data;                                                                                 // cmd_xbar_demux:src14_data -> burst_adapter_014:sink0_data
	wire   [18:0] cmd_xbar_demux_src14_channel;                                                                              // cmd_xbar_demux:src14_channel -> burst_adapter_014:sink0_channel
	wire          cmd_xbar_demux_src16_endofpacket;                                                                          // cmd_xbar_demux:src16_endofpacket -> burst_adapter_016:sink0_endofpacket
	wire          cmd_xbar_demux_src16_valid;                                                                                // cmd_xbar_demux:src16_valid -> burst_adapter_016:sink0_valid
	wire          cmd_xbar_demux_src16_startofpacket;                                                                        // cmd_xbar_demux:src16_startofpacket -> burst_adapter_016:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src16_data;                                                                                 // cmd_xbar_demux:src16_data -> burst_adapter_016:sink0_data
	wire   [18:0] cmd_xbar_demux_src16_channel;                                                                              // cmd_xbar_demux:src16_channel -> burst_adapter_016:sink0_channel
	wire          cmd_xbar_demux_src17_endofpacket;                                                                          // cmd_xbar_demux:src17_endofpacket -> burst_adapter_017:sink0_endofpacket
	wire          cmd_xbar_demux_src17_valid;                                                                                // cmd_xbar_demux:src17_valid -> burst_adapter_017:sink0_valid
	wire          cmd_xbar_demux_src17_startofpacket;                                                                        // cmd_xbar_demux:src17_startofpacket -> burst_adapter_017:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src17_data;                                                                                 // cmd_xbar_demux:src17_data -> burst_adapter_017:sink0_data
	wire   [18:0] cmd_xbar_demux_src17_channel;                                                                              // cmd_xbar_demux:src17_channel -> burst_adapter_017:sink0_channel
	wire          cmd_xbar_demux_src18_endofpacket;                                                                          // cmd_xbar_demux:src18_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	wire          cmd_xbar_demux_src18_valid;                                                                                // cmd_xbar_demux:src18_valid -> cmd_xbar_mux_018:sink0_valid
	wire          cmd_xbar_demux_src18_startofpacket;                                                                        // cmd_xbar_demux:src18_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src18_data;                                                                                 // cmd_xbar_demux:src18_data -> cmd_xbar_mux_018:sink0_data
	wire   [18:0] cmd_xbar_demux_src18_channel;                                                                              // cmd_xbar_demux:src18_channel -> cmd_xbar_mux_018:sink0_channel
	wire          cmd_xbar_demux_src18_ready;                                                                                // cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux:src18_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                       // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                             // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                     // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src0_data;                                                                              // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src0_channel;                                                                           // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                             // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                       // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                             // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                     // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src1_data;                                                                              // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_002:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src1_channel;                                                                           // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                             // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                       // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                             // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                     // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src2_data;                                                                              // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_005:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src2_channel;                                                                           // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                             // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                       // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                             // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_006:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                     // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src3_data;                                                                              // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_006:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src3_channel;                                                                           // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                             // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                       // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                             // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_018:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                     // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src4_data;                                                                              // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_018:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src4_channel;                                                                           // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_018:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                             // cmd_xbar_mux_018:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                           // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                 // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                         // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [107:0] rsp_xbar_demux_src0_data;                                                                                  // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [18:0] rsp_xbar_demux_src0_channel;                                                                               // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                 // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                           // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                 // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                         // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [107:0] rsp_xbar_demux_src1_data;                                                                                  // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [18:0] rsp_xbar_demux_src1_channel;                                                                               // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                 // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                       // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                             // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                     // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [107:0] rsp_xbar_demux_001_src0_data;                                                                              // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [18:0] rsp_xbar_demux_001_src0_channel;                                                                           // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                             // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                       // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                             // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                     // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [107:0] rsp_xbar_demux_002_src0_data;                                                                              // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [18:0] rsp_xbar_demux_002_src0_channel;                                                                           // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                             // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                       // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                             // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                     // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [107:0] rsp_xbar_demux_002_src1_data;                                                                              // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [18:0] rsp_xbar_demux_002_src1_channel;                                                                           // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                             // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                       // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                             // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                     // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [107:0] rsp_xbar_demux_003_src0_data;                                                                              // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [18:0] rsp_xbar_demux_003_src0_channel;                                                                           // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                             // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                       // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                             // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                     // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [107:0] rsp_xbar_demux_004_src0_data;                                                                              // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src0_channel;                                                                           // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                             // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                       // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                             // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                     // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [107:0] rsp_xbar_demux_005_src0_data;                                                                              // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src0_channel;                                                                           // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                             // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                       // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                             // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                     // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [107:0] rsp_xbar_demux_005_src1_data;                                                                              // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [18:0] rsp_xbar_demux_005_src1_channel;                                                                           // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                             // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                       // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                             // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                     // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [107:0] rsp_xbar_demux_006_src0_data;                                                                              // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [18:0] rsp_xbar_demux_006_src0_channel;                                                                           // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                             // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                                       // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                             // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                                     // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [107:0] rsp_xbar_demux_006_src1_data;                                                                              // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [18:0] rsp_xbar_demux_006_src1_channel;                                                                           // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                             // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_006:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                       // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                             // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                     // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [107:0] rsp_xbar_demux_007_src0_data;                                                                              // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src0_channel;                                                                           // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                             // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                       // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                             // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                     // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [107:0] rsp_xbar_demux_008_src0_data;                                                                              // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire   [18:0] rsp_xbar_demux_008_src0_channel;                                                                           // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                             // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                       // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                             // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                     // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [107:0] rsp_xbar_demux_009_src0_data;                                                                              // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src0_channel;                                                                           // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                             // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                       // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                             // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                     // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [107:0] rsp_xbar_demux_010_src0_data;                                                                              // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src0_channel;                                                                           // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                             // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                       // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                             // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                     // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [107:0] rsp_xbar_demux_011_src0_data;                                                                              // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire   [18:0] rsp_xbar_demux_011_src0_channel;                                                                           // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                             // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                       // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                             // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                     // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [107:0] rsp_xbar_demux_012_src0_data;                                                                              // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire   [18:0] rsp_xbar_demux_012_src0_channel;                                                                           // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                             // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                       // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                             // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                     // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [107:0] rsp_xbar_demux_013_src0_data;                                                                              // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire   [18:0] rsp_xbar_demux_013_src0_channel;                                                                           // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                             // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                       // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                             // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                     // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [107:0] rsp_xbar_demux_014_src0_data;                                                                              // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire   [18:0] rsp_xbar_demux_014_src0_channel;                                                                           // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                             // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                       // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                             // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                     // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [107:0] rsp_xbar_demux_016_src0_data;                                                                              // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire   [18:0] rsp_xbar_demux_016_src0_channel;                                                                           // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                             // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                       // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                             // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                     // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [107:0] rsp_xbar_demux_017_src0_data;                                                                              // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire   [18:0] rsp_xbar_demux_017_src0_channel;                                                                           // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                             // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                       // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                             // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                     // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	wire  [107:0] rsp_xbar_demux_018_src0_data;                                                                              // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux:sink18_data
	wire   [18:0] rsp_xbar_demux_018_src0_channel;                                                                           // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                             // rsp_xbar_mux:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_018_src1_endofpacket;                                                                       // rsp_xbar_demux_018:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_018_src1_valid;                                                                             // rsp_xbar_demux_018:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_018_src1_startofpacket;                                                                     // rsp_xbar_demux_018:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [107:0] rsp_xbar_demux_018_src1_data;                                                                              // rsp_xbar_demux_018:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [18:0] rsp_xbar_demux_018_src1_channel;                                                                           // rsp_xbar_demux_018:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_018_src1_ready;                                                                             // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_018:src1_ready
	wire          limiter_cmd_src_endofpacket;                                                                               // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                             // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [107:0] limiter_cmd_src_data;                                                                                      // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [18:0] limiter_cmd_src_channel;                                                                                   // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                     // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                              // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                    // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                            // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [107:0] rsp_xbar_mux_src_data;                                                                                     // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_src_channel;                                                                                  // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                    // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                           // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                         // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [107:0] limiter_001_cmd_src_data;                                                                                  // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [18:0] limiter_001_cmd_src_channel;                                                                               // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                 // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                          // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                        // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [107:0] rsp_xbar_mux_001_src_data;                                                                                 // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_001_src_channel;                                                                              // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                              // cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                    // cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                            // cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [107:0] cmd_xbar_mux_src_data;                                                                                     // cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	wire   [18:0] cmd_xbar_mux_src_channel;                                                                                  // cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_src_ready;                                                                                    // burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                 // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                       // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                               // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [107:0] id_router_src_data;                                                                                        // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [18:0] id_router_src_channel;                                                                                     // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                       // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                                                 // burst_adapter_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                                             // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                   // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                           // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [107:0] id_router_003_src_data;                                                                                    // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [18:0] id_router_003_src_channel;                                                                                 // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                   // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_src4_ready;                                                                                 // burst_adapter_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          id_router_004_src_endofpacket;                                                                             // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                   // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                           // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [107:0] id_router_004_src_data;                                                                                    // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [18:0] id_router_004_src_channel;                                                                                 // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                   // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                          // cmd_xbar_mux_005:src_endofpacket -> burst_adapter_005:sink0_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                // cmd_xbar_mux_005:src_valid -> burst_adapter_005:sink0_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                        // cmd_xbar_mux_005:src_startofpacket -> burst_adapter_005:sink0_startofpacket
	wire  [107:0] cmd_xbar_mux_005_src_data;                                                                                 // cmd_xbar_mux_005:src_data -> burst_adapter_005:sink0_data
	wire   [18:0] cmd_xbar_mux_005_src_channel;                                                                              // cmd_xbar_mux_005:src_channel -> burst_adapter_005:sink0_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                // burst_adapter_005:sink0_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                             // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                   // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                           // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [107:0] id_router_005_src_data;                                                                                    // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [18:0] id_router_005_src_channel;                                                                                 // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                   // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_src7_ready;                                                                                 // burst_adapter_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire          id_router_007_src_endofpacket;                                                                             // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                   // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                           // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [107:0] id_router_007_src_data;                                                                                    // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [18:0] id_router_007_src_channel;                                                                                 // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                   // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_src8_ready;                                                                                 // burst_adapter_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire          id_router_008_src_endofpacket;                                                                             // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                   // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                           // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [107:0] id_router_008_src_data;                                                                                    // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [18:0] id_router_008_src_channel;                                                                                 // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                   // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_src9_ready;                                                                                 // burst_adapter_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire          id_router_009_src_endofpacket;                                                                             // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                   // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                           // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [107:0] id_router_009_src_data;                                                                                    // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [18:0] id_router_009_src_channel;                                                                                 // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                   // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_src10_ready;                                                                                // burst_adapter_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire          id_router_010_src_endofpacket;                                                                             // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                   // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                           // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [107:0] id_router_010_src_data;                                                                                    // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [18:0] id_router_010_src_channel;                                                                                 // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                   // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_src11_ready;                                                                                // burst_adapter_011:sink0_ready -> cmd_xbar_demux:src11_ready
	wire          id_router_011_src_endofpacket;                                                                             // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                   // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                           // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [107:0] id_router_011_src_data;                                                                                    // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [18:0] id_router_011_src_channel;                                                                                 // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                   // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_src12_ready;                                                                                // burst_adapter_012:sink0_ready -> cmd_xbar_demux:src12_ready
	wire          id_router_012_src_endofpacket;                                                                             // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                   // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                           // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [107:0] id_router_012_src_data;                                                                                    // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [18:0] id_router_012_src_channel;                                                                                 // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                   // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_src13_ready;                                                                                // burst_adapter_013:sink0_ready -> cmd_xbar_demux:src13_ready
	wire          id_router_013_src_endofpacket;                                                                             // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                   // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                           // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [107:0] id_router_013_src_data;                                                                                    // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [18:0] id_router_013_src_channel;                                                                                 // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                   // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_src14_ready;                                                                                // burst_adapter_014:sink0_ready -> cmd_xbar_demux:src14_ready
	wire          id_router_014_src_endofpacket;                                                                             // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                   // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                           // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [107:0] id_router_014_src_data;                                                                                    // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [18:0] id_router_014_src_channel;                                                                                 // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                   // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          crosser_out_ready;                                                                                         // burst_adapter_015:sink0_ready -> crosser:out_ready
	wire          id_router_015_src_endofpacket;                                                                             // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                   // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                           // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [107:0] id_router_015_src_data;                                                                                    // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [18:0] id_router_015_src_channel;                                                                                 // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                   // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_src16_ready;                                                                                // burst_adapter_016:sink0_ready -> cmd_xbar_demux:src16_ready
	wire          id_router_016_src_endofpacket;                                                                             // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                   // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                           // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [107:0] id_router_016_src_data;                                                                                    // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [18:0] id_router_016_src_channel;                                                                                 // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                   // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_src17_ready;                                                                                // burst_adapter_017:sink0_ready -> cmd_xbar_demux:src17_ready
	wire          id_router_017_src_endofpacket;                                                                             // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                   // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                           // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [107:0] id_router_017_src_data;                                                                                    // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [18:0] id_router_017_src_channel;                                                                                 // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                   // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_src1_ready;                                                                                 // width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_src_endofpacket;                                                                             // width_adapter:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                   // width_adapter:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                           // width_adapter:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [80:0] width_adapter_src_data;                                                                                    // width_adapter:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_src_ready;                                                                                   // burst_adapter_001:sink0_ready -> width_adapter:out_ready
	wire   [18:0] width_adapter_src_channel;                                                                                 // width_adapter:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                             // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                                   // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                           // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [80:0] id_router_001_src_data;                                                                                    // id_router_001:src_data -> width_adapter_001:in_data
	wire   [18:0] id_router_001_src_channel;                                                                                 // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                                   // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                         // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                               // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                       // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [107:0] width_adapter_001_src_data;                                                                                // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                               // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [18:0] width_adapter_001_src_channel;                                                                             // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                          // cmd_xbar_mux_002:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                // cmd_xbar_mux_002:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                        // cmd_xbar_mux_002:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [107:0] cmd_xbar_mux_002_src_data;                                                                                 // cmd_xbar_mux_002:src_data -> width_adapter_002:in_data
	wire   [18:0] cmd_xbar_mux_002_src_channel;                                                                              // cmd_xbar_mux_002:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                // width_adapter_002:in_ready -> cmd_xbar_mux_002:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                         // width_adapter_002:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                               // width_adapter_002:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                       // width_adapter_002:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [89:0] width_adapter_002_src_data;                                                                                // width_adapter_002:out_data -> burst_adapter_002:sink0_data
	wire          width_adapter_002_src_ready;                                                                               // burst_adapter_002:sink0_ready -> width_adapter_002:out_ready
	wire   [18:0] width_adapter_002_src_channel;                                                                             // width_adapter_002:out_channel -> burst_adapter_002:sink0_channel
	wire          id_router_002_src_endofpacket;                                                                             // id_router_002:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_002_src_valid;                                                                                   // id_router_002:src_valid -> width_adapter_003:in_valid
	wire          id_router_002_src_startofpacket;                                                                           // id_router_002:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [89:0] id_router_002_src_data;                                                                                    // id_router_002:src_data -> width_adapter_003:in_data
	wire   [18:0] id_router_002_src_channel;                                                                                 // id_router_002:src_channel -> width_adapter_003:in_channel
	wire          id_router_002_src_ready;                                                                                   // width_adapter_003:in_ready -> id_router_002:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                         // width_adapter_003:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                               // width_adapter_003:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                       // width_adapter_003:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [107:0] width_adapter_003_src_data;                                                                                // width_adapter_003:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_003_src_ready;                                                                               // rsp_xbar_demux_002:sink_ready -> width_adapter_003:out_ready
	wire   [18:0] width_adapter_003_src_channel;                                                                             // width_adapter_003:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                          // cmd_xbar_mux_006:src_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                                // cmd_xbar_mux_006:src_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                                        // cmd_xbar_mux_006:src_startofpacket -> width_adapter_004:in_startofpacket
	wire  [107:0] cmd_xbar_mux_006_src_data;                                                                                 // cmd_xbar_mux_006:src_data -> width_adapter_004:in_data
	wire   [18:0] cmd_xbar_mux_006_src_channel;                                                                              // cmd_xbar_mux_006:src_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                                // width_adapter_004:in_ready -> cmd_xbar_mux_006:src_ready
	wire          width_adapter_004_src_endofpacket;                                                                         // width_adapter_004:out_endofpacket -> burst_adapter_006:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                               // width_adapter_004:out_valid -> burst_adapter_006:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                       // width_adapter_004:out_startofpacket -> burst_adapter_006:sink0_startofpacket
	wire   [89:0] width_adapter_004_src_data;                                                                                // width_adapter_004:out_data -> burst_adapter_006:sink0_data
	wire          width_adapter_004_src_ready;                                                                               // burst_adapter_006:sink0_ready -> width_adapter_004:out_ready
	wire   [18:0] width_adapter_004_src_channel;                                                                             // width_adapter_004:out_channel -> burst_adapter_006:sink0_channel
	wire          id_router_006_src_endofpacket;                                                                             // id_router_006:src_endofpacket -> width_adapter_005:in_endofpacket
	wire          id_router_006_src_valid;                                                                                   // id_router_006:src_valid -> width_adapter_005:in_valid
	wire          id_router_006_src_startofpacket;                                                                           // id_router_006:src_startofpacket -> width_adapter_005:in_startofpacket
	wire   [89:0] id_router_006_src_data;                                                                                    // id_router_006:src_data -> width_adapter_005:in_data
	wire   [18:0] id_router_006_src_channel;                                                                                 // id_router_006:src_channel -> width_adapter_005:in_channel
	wire          id_router_006_src_ready;                                                                                   // width_adapter_005:in_ready -> id_router_006:src_ready
	wire          width_adapter_005_src_endofpacket;                                                                         // width_adapter_005:out_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          width_adapter_005_src_valid;                                                                               // width_adapter_005:out_valid -> rsp_xbar_demux_006:sink_valid
	wire          width_adapter_005_src_startofpacket;                                                                       // width_adapter_005:out_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [107:0] width_adapter_005_src_data;                                                                                // width_adapter_005:out_data -> rsp_xbar_demux_006:sink_data
	wire          width_adapter_005_src_ready;                                                                               // rsp_xbar_demux_006:sink_ready -> width_adapter_005:out_ready
	wire   [18:0] width_adapter_005_src_channel;                                                                             // width_adapter_005:out_channel -> rsp_xbar_demux_006:sink_channel
	wire          cmd_xbar_mux_018_src_endofpacket;                                                                          // cmd_xbar_mux_018:src_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_mux_018_src_valid;                                                                                // cmd_xbar_mux_018:src_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_mux_018_src_startofpacket;                                                                        // cmd_xbar_mux_018:src_startofpacket -> width_adapter_006:in_startofpacket
	wire  [107:0] cmd_xbar_mux_018_src_data;                                                                                 // cmd_xbar_mux_018:src_data -> width_adapter_006:in_data
	wire   [18:0] cmd_xbar_mux_018_src_channel;                                                                              // cmd_xbar_mux_018:src_channel -> width_adapter_006:in_channel
	wire          cmd_xbar_mux_018_src_ready;                                                                                // width_adapter_006:in_ready -> cmd_xbar_mux_018:src_ready
	wire          width_adapter_006_src_endofpacket;                                                                         // width_adapter_006:out_endofpacket -> burst_adapter_018:sink0_endofpacket
	wire          width_adapter_006_src_valid;                                                                               // width_adapter_006:out_valid -> burst_adapter_018:sink0_valid
	wire          width_adapter_006_src_startofpacket;                                                                       // width_adapter_006:out_startofpacket -> burst_adapter_018:sink0_startofpacket
	wire   [80:0] width_adapter_006_src_data;                                                                                // width_adapter_006:out_data -> burst_adapter_018:sink0_data
	wire          width_adapter_006_src_ready;                                                                               // burst_adapter_018:sink0_ready -> width_adapter_006:out_ready
	wire   [18:0] width_adapter_006_src_channel;                                                                             // width_adapter_006:out_channel -> burst_adapter_018:sink0_channel
	wire          id_router_018_src_endofpacket;                                                                             // id_router_018:src_endofpacket -> width_adapter_007:in_endofpacket
	wire          id_router_018_src_valid;                                                                                   // id_router_018:src_valid -> width_adapter_007:in_valid
	wire          id_router_018_src_startofpacket;                                                                           // id_router_018:src_startofpacket -> width_adapter_007:in_startofpacket
	wire   [80:0] id_router_018_src_data;                                                                                    // id_router_018:src_data -> width_adapter_007:in_data
	wire   [18:0] id_router_018_src_channel;                                                                                 // id_router_018:src_channel -> width_adapter_007:in_channel
	wire          id_router_018_src_ready;                                                                                   // width_adapter_007:in_ready -> id_router_018:src_ready
	wire          width_adapter_007_src_endofpacket;                                                                         // width_adapter_007:out_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          width_adapter_007_src_valid;                                                                               // width_adapter_007:out_valid -> rsp_xbar_demux_018:sink_valid
	wire          width_adapter_007_src_startofpacket;                                                                       // width_adapter_007:out_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [107:0] width_adapter_007_src_data;                                                                                // width_adapter_007:out_data -> rsp_xbar_demux_018:sink_data
	wire          width_adapter_007_src_ready;                                                                               // rsp_xbar_demux_018:sink_ready -> width_adapter_007:out_ready
	wire   [18:0] width_adapter_007_src_channel;                                                                             // width_adapter_007:out_channel -> rsp_xbar_demux_018:sink_channel
	wire          crosser_out_endofpacket;                                                                                   // crosser:out_endofpacket -> burst_adapter_015:sink0_endofpacket
	wire          crosser_out_valid;                                                                                         // crosser:out_valid -> burst_adapter_015:sink0_valid
	wire          crosser_out_startofpacket;                                                                                 // crosser:out_startofpacket -> burst_adapter_015:sink0_startofpacket
	wire  [107:0] crosser_out_data;                                                                                          // crosser:out_data -> burst_adapter_015:sink0_data
	wire   [18:0] crosser_out_channel;                                                                                       // crosser:out_channel -> burst_adapter_015:sink0_channel
	wire          cmd_xbar_demux_src15_endofpacket;                                                                          // cmd_xbar_demux:src15_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src15_valid;                                                                                // cmd_xbar_demux:src15_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src15_startofpacket;                                                                        // cmd_xbar_demux:src15_startofpacket -> crosser:in_startofpacket
	wire  [107:0] cmd_xbar_demux_src15_data;                                                                                 // cmd_xbar_demux:src15_data -> crosser:in_data
	wire   [18:0] cmd_xbar_demux_src15_channel;                                                                              // cmd_xbar_demux:src15_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src15_ready;                                                                                // crosser:in_ready -> cmd_xbar_demux:src15_ready
	wire          crosser_001_out_endofpacket;                                                                               // crosser_001:out_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire          crosser_001_out_valid;                                                                                     // crosser_001:out_valid -> rsp_xbar_mux:sink15_valid
	wire          crosser_001_out_startofpacket;                                                                             // crosser_001:out_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [107:0] crosser_001_out_data;                                                                                      // crosser_001:out_data -> rsp_xbar_mux:sink15_data
	wire   [18:0] crosser_001_out_channel;                                                                                   // crosser_001:out_channel -> rsp_xbar_mux:sink15_channel
	wire          crosser_001_out_ready;                                                                                     // rsp_xbar_mux:sink15_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                       // rsp_xbar_demux_015:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                             // rsp_xbar_demux_015:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                     // rsp_xbar_demux_015:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [107:0] rsp_xbar_demux_015_src0_data;                                                                              // rsp_xbar_demux_015:src0_data -> crosser_001:in_data
	wire   [18:0] rsp_xbar_demux_015_src0_channel;                                                                           // rsp_xbar_demux_015:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                             // crosser_001:in_ready -> rsp_xbar_demux_015:src0_ready
	wire   [18:0] limiter_cmd_valid_data;                                                                                    // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [18:0] limiter_001_cmd_valid_data;                                                                                // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                  // timer:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                  // add_button:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                  // remove_button:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                  // cancel_button:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                  // switch:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                                  // barcode_scanner_ps2:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver8_irq;                                                                                  // dm9000a_if_ethernet:avs_s1_irq_oINT -> irq_mapper:receiver8_irq
	wire   [31:0] nios2_qsys_d_irq_irq;                                                                                      // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire          irq_mapper_receiver7_irq;                                                                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver7_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                             // audio_core:irq -> irq_synchronizer:receiver_irq

	niosII_system_nios2_qsys nios2_qsys (
		.clk                                   (main_pll_sys_clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.d_burstcount                          (nios2_qsys_data_master_burstcount),                                         //                          .burstcount
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_burstcount                          (nios2_qsys_instruction_master_burstcount),                                  //                          .burstcount
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	niosII_system_onchip_memory2 onchip_memory2 (
		.clk        (main_pll_sys_clk_clk),                                        //   clk1.clk
		.address    (onchip_memory2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                               // reset1.reset
	);

	niosII_system_sysid_qsys sysid_qsys (
		.clock    (main_pll_sys_clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.readdata (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	niosII_system_timer timer (
		.clk        (main_pll_sys_clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                            //   irq.irq
	);

	niosII_system_jtag_uart jtag_uart (
		.clk            (main_pll_sys_clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	niosII_system_character_lcd character_lcd (
		.clk         (main_pll_sys_clk_clk),                                                      //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                            //  clock_reset_reset.reset
		.address     (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (character_lcd_external_interface_DATA),                                     // external_interface.export
		.LCD_ON      (character_lcd_external_interface_ON),                                       //                   .export
		.LCD_BLON    (character_lcd_external_interface_BLON),                                     //                   .export
		.LCD_EN      (character_lcd_external_interface_EN),                                       //                   .export
		.LCD_RS      (character_lcd_external_interface_RS),                                       //                   .export
		.LCD_RW      (character_lcd_external_interface_RW)                                        //                   .export
	);

	niosII_system_green_leds green_leds (
		.clk        (main_pll_sys_clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (green_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~green_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (green_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (green_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (green_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (green_leds_external_connection_export)                    // external_connection.export
	);

	niosII_system_switch switch (
		.clk        (main_pll_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (switch_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                             //                 irq.irq
	);

	niosII_system_sdram sdram (
		.clk            (main_pll_sys_clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	niosII_system_sram sram (
		.clk           (main_pll_sys_clk_clk),                                                //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                      //  clock_reset_reset.reset
		.SRAM_DQ       (sram_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_external_interface_WE_N),                                        //                   .export
		.address       (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	niosII_system_add_button add_button (
		.clk        (main_pll_sys_clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (add_button_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~add_button_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (add_button_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (add_button_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (add_button_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (add_button_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                                 //                 irq.irq
	);

	niosII_system_add_button remove_button (
		.clk        (main_pll_sys_clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (remove_button_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~remove_button_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (remove_button_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (remove_button_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (remove_button_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (remove_button_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                                    //                 irq.irq
	);

	niosII_system_add_button cancel_button (
		.clk        (main_pll_sys_clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (cancel_button_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~cancel_button_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (cancel_button_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (cancel_button_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (cancel_button_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (cancel_button_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                                    //                 irq.irq
	);

	niosII_system_green_leds red_leds (
		.clk        (main_pll_sys_clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (red_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~red_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (red_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (red_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (red_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (red_leds_external_connection_export)                    // external_connection.export
	);

	niosII_system_barcode_scanner_ps2 barcode_scanner_ps2 (
		.clk         (main_pll_sys_clk_clk),                                                            //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                                  //  clock_reset_reset.reset
		.address     (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_address),     //   avalon_ps2_slave.address
		.chipselect  (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.byteenable  (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.read        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver6_irq),                                                        //          interrupt.irq
		.PS2_CLK     (barcode_scanner_ps2_external_interface_CLK),                                      // external_interface.export
		.PS2_DAT     (barcode_scanner_ps2_external_interface_DAT)                                       //                   .export
	);

	niosII_system_audio_core audio_core (
		.clk         (main_pll_audio_clk_clk),                                                  //        clock_reset.clk
		.reset       (rst_controller_001_reset_out_reset),                                      //  clock_reset_reset.reset
		.address     (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_address),    // avalon_audio_slave.address
		.chipselect  (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read        (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write       (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata   (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata    (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq         (irq_synchronizer_receiver_irq),                                           //          interrupt.irq
		.AUD_ADCDAT  (audio_core_external_interface_ADCDAT),                                    // external_interface.export
		.AUD_ADCLRCK (audio_core_external_interface_ADCLRCK),                                   //                   .export
		.AUD_BCLK    (audio_core_external_interface_BCLK),                                      //                   .export
		.AUD_DACDAT  (audio_core_external_interface_DACDAT),                                    //                   .export
		.AUD_DACLRCK (audio_core_external_interface_DACLRCK)                                    //                   .export
	);

	niosII_system_audio_config audio_config (
		.clk         (main_pll_sys_clk_clk),                                                           //            clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                                 //      clock_reset_reset.reset
		.address     (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_config_external_interface_SDAT),                                           //     external_interface.export
		.I2C_SCLK    (audio_config_external_interface_SCLK)                                            //                       .export
	);

	niosII_system_main_pll main_pll (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_002_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (main_pll_sys_clk_clk),               //              sys_clk.clk
		.sys_reset_n (main_pll_sys_clk_reset_reset),       //        sys_clk_reset.reset_n
		.SDRAM_CLK   (main_pll_sdram_clk_clk),             //            sdram_clk.clk
		.CLOCK_27    (clock_27mhz_clk_in_clk),             //     clk_in_secondary.clk
		.AUD_CLK     (main_pll_audio_clk_clk)              //            audio_clk.clk
	);

	DM9000A_IF dm9000a_if_ethernet (
		.avs_s1_clk_iCLK           (main_pll_sys_clk_clk),                                              //       s1_clock.clk
		.avs_s1_reset_n_iRST_N     (~rst_controller_reset_out_reset),                                   // s1_clock_reset.reset_n
		.avs_s1_writedata_iDATA    (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_writedata),   //             s1.writedata
		.avs_s1_readdata_oDATA     (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.avs_s1_address_iCMD       (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_address),     //               .address
		.avs_s1_read_n_iRD_N       (~dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_read),       //               .read_n
		.avs_s1_write_n_iWR_N      (~dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_write),      //               .write_n
		.avs_s1_chipselect_n_iCS_N (~dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.avs_s1_irq_oINT           (irq_mapper_receiver8_irq),                                          //         s1_irq.irq
		.avs_s1_export_ENET_DATA   (dm9000a_if_ethernet_s1_export_DATA),                                //      s1_export.export
		.avs_s1_export_ENET_CMD    (dm9000a_if_ethernet_s1_export_CMD),                                 //               .export
		.avs_s1_export_ENET_RD_N   (dm9000a_if_ethernet_s1_export_RD_N),                                //               .export
		.avs_s1_export_ENET_WR_N   (dm9000a_if_ethernet_s1_export_WR_N),                                //               .export
		.avs_s1_export_ENET_CS_N   (dm9000a_if_ethernet_s1_export_CS_N),                                //               .export
		.avs_s1_export_ENET_RST_N  (dm9000a_if_ethernet_s1_export_RST_N),                               //               .export
		.avs_s1_export_ENET_INT    (dm9000a_if_ethernet_s1_export_INT),                                 //               .export
		.avs_s1_export_ENET_CLK    (dm9000a_if_ethernet_s1_export_CLK)                                  //               .export
	);

	niosII_system_tristate_controller #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) tristate_controller (
		.clk_clk               (main_pll_sys_clk_clk),                                                 //   clk.clk
		.reset_reset           (rst_controller_reset_out_reset),                                       // reset.reset
		.uas_address           (tristate_controller_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount        (tristate_controller_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read              (tristate_controller_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write             (tristate_controller_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest       (tristate_controller_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid     (tristate_controller_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable        (tristate_controller_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata          (tristate_controller_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata         (tristate_controller_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock              (tristate_controller_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess       (tristate_controller_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out       (tristate_controller_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out        (tristate_controller_tcm_read_n_out),                                   //      .read_n_out
		.tcm_begintransfer_out (tristate_controller_tcm_begintransfer_out),                            //      .begintransfer_out
		.tcm_chipselect_n_out  (tristate_controller_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request           (tristate_controller_tcm_request),                                      //      .request
		.tcm_grant             (tristate_controller_tcm_grant),                                        //      .grant
		.tcm_address_out       (tristate_controller_tcm_address_out),                                  //      .address_out
		.tcm_byteenable_out    (tristate_controller_tcm_byteenable_out),                               //      .byteenable_out
		.tcm_data_out          (tristate_controller_tcm_data_out),                                     //      .data_out
		.tcm_data_outen        (tristate_controller_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in           (tristate_controller_tcm_data_in)                                       //      .data_in
	);

	niosII_system_tristate_conduit_bridge tristate_conduit_bridge (
		.clk                                           (main_pll_sys_clk_clk),                                                          //   clk.clk
		.reset                                         (rst_controller_reset_out_reset),                                                // reset.reset
		.request                                       (tristate_conduit_pin_sharer_tcm_request),                                       //   tcs.request
		.grant                                         (tristate_conduit_pin_sharer_tcm_grant),                                         //      .grant
		.tcs_tristate_controller_tcm_read_n_out        (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_read_n_out_out),        //      .tristate_controller_tcm_read_n_out_out
		.tcs_tristate_controller_tcm_address_out       (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_address_out_out),       //      .tristate_controller_tcm_address_out_out
		.tcs_tristate_controller_tcm_data_out          (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_out),          //      .tristate_controller_tcm_data_out_out
		.tcs_tristate_controller_tcm_data_outen        (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_outen),        //      .tristate_controller_tcm_data_out_outen
		.tcs_tristate_controller_tcm_data_in           (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_in),           //      .tristate_controller_tcm_data_out_in
		.tcs_tristate_controller_tcm_byteenable_out    (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_byteenable_out_out),    //      .tristate_controller_tcm_byteenable_out_out
		.tcs_tristate_controller_tcm_begintransfer_out (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_begintransfer_out_out), //      .tristate_controller_tcm_begintransfer_out_out
		.tcs_tristate_controller_tcm_write_n_out       (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_write_n_out_out),       //      .tristate_controller_tcm_write_n_out_out
		.tcs_tristate_controller_tcm_chipselect_n_out  (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_chipselect_n_out_out),  //      .tristate_controller_tcm_chipselect_n_out_out
		.tristate_controller_tcm_read_n_out            (tristate_conduit_bridge_out_tristate_controller_tcm_read_n_out),                //   out.tristate_controller_tcm_read_n_out
		.tristate_controller_tcm_address_out           (tristate_conduit_bridge_out_tristate_controller_tcm_address_out),               //      .tristate_controller_tcm_address_out
		.tristate_controller_tcm_data_out              (tristate_conduit_bridge_out_tristate_controller_tcm_data_out),                  //      .tristate_controller_tcm_data_out
		.tristate_controller_tcm_byteenable_out        (tristate_conduit_bridge_out_tristate_controller_tcm_byteenable_out),            //      .tristate_controller_tcm_byteenable_out
		.tristate_controller_tcm_begintransfer_out     (tristate_conduit_bridge_out_tristate_controller_tcm_begintransfer_out),         //      .tristate_controller_tcm_begintransfer_out
		.tristate_controller_tcm_write_n_out           (tristate_conduit_bridge_out_tristate_controller_tcm_write_n_out),               //      .tristate_controller_tcm_write_n_out
		.tristate_controller_tcm_chipselect_n_out      (tristate_conduit_bridge_out_tristate_controller_tcm_chipselect_n_out)           //      .tristate_controller_tcm_chipselect_n_out
	);

	niosII_system_tristate_conduit_pin_sharer tristate_conduit_pin_sharer (
		.clk_clk                                   (main_pll_sys_clk_clk),                                                          //   clk.clk
		.reset_reset                               (rst_controller_reset_out_reset),                                                // reset.reset
		.request                                   (tristate_conduit_pin_sharer_tcm_request),                                       //   tcm.request
		.grant                                     (tristate_conduit_pin_sharer_tcm_grant),                                         //      .grant
		.tristate_controller_tcm_byteenable_out    (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_byteenable_out_out),    //      .tristate_controller_tcm_byteenable_out_out
		.tristate_controller_tcm_address_out       (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_address_out_out),       //      .tristate_controller_tcm_address_out_out
		.tristate_controller_tcm_read_n_out        (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_read_n_out_out),        //      .tristate_controller_tcm_read_n_out_out
		.tristate_controller_tcm_write_n_out       (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_write_n_out_out),       //      .tristate_controller_tcm_write_n_out_out
		.tristate_controller_tcm_data_out          (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_out),          //      .tristate_controller_tcm_data_out_out
		.tristate_controller_tcm_data_in           (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_in),           //      .tristate_controller_tcm_data_out_in
		.tristate_controller_tcm_data_outen        (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_data_out_outen),        //      .tristate_controller_tcm_data_out_outen
		.tristate_controller_tcm_chipselect_n_out  (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_chipselect_n_out_out),  //      .tristate_controller_tcm_chipselect_n_out_out
		.tristate_controller_tcm_begintransfer_out (tristate_conduit_pin_sharer_tcm_tristate_controller_tcm_begintransfer_out_out), //      .tristate_controller_tcm_begintransfer_out_out
		.tcs0_request                              (tristate_controller_tcm_request),                                               //  tcs0.request
		.tcs0_grant                                (tristate_controller_tcm_grant),                                                 //      .grant
		.tcs0_byteenable_out                       (tristate_controller_tcm_byteenable_out),                                        //      .byteenable_out
		.tcs0_address_out                          (tristate_controller_tcm_address_out),                                           //      .address_out
		.tcs0_read_n_out                           (tristate_controller_tcm_read_n_out),                                            //      .read_n_out
		.tcs0_write_n_out                          (tristate_controller_tcm_write_n_out),                                           //      .write_n_out
		.tcs0_data_out                             (tristate_controller_tcm_data_out),                                              //      .data_out
		.tcs0_data_in                              (tristate_controller_tcm_data_in),                                               //      .data_in
		.tcs0_data_outen                           (tristate_controller_tcm_data_outen),                                            //      .data_outen
		.tcs0_chipselect_n_out                     (tristate_controller_tcm_chipselect_n_out),                                      //      .chipselect_n_out
		.tcs0_begintransfer_out                    (tristate_controller_tcm_begintransfer_out)                                      //      .begintransfer_out
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_data_master_translator (
		.clk                   (main_pll_sys_clk_clk),                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (nios2_qsys_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (nios2_qsys_data_master_burstcount),                                         //                          .burstcount
		.av_byteenable         (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_qsys_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_instruction_master_translator (
		.clk                   (main_pll_sys_clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (nios2_qsys_instruction_master_burstcount),                                         //                          .burstcount
		.av_read               (nios2_qsys_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable         (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_write              (1'b0),                                                                             //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_jtag_debug_module_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_avalon_lcd_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (character_lcd_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_byteenable         (),                                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_debugaccess        (),                                                                                          //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_avalon_sram_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_control_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                    //              (terminated)
		.av_read               (),                                                                                    //              (terminated)
		.av_writedata          (),                                                                                    //              (terminated)
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (green_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (green_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (green_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (green_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (green_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (switch_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (switch_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (switch_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (switch_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) add_button_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (add_button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (add_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (add_button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (add_button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (add_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (add_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (add_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (add_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (add_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (add_button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (add_button_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (add_button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (add_button_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (add_button_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) remove_button_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (remove_button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (remove_button_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (remove_button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (remove_button_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (remove_button_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cancel_button_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cancel_button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cancel_button_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cancel_button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cancel_button_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (cancel_button_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) red_leds_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (red_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (red_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (red_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (red_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (red_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) barcode_scanner_ps2_avalon_ps2_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                                //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_core_avalon_audio_slave_translator (
		.clk                   (main_pll_audio_clk_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (audio_core_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_config_avalon_av_config_slave_translator (
		.clk                   (main_pll_sys_clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                 //                    reset.reset
		.uav_address           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (audio_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                               //              (terminated)
		.av_lock               (),                                                                                               //              (terminated)
		.av_chipselect         (),                                                                                               //              (terminated)
		.av_clken              (),                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (3),
		.AV_WRITE_WAIT_CYCLES           (3),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (1)
	) dm9000a_if_ethernet_s1_translator (
		.clk                   (main_pll_sys_clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (dm9000a_if_ethernet_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tristate_controller_uas_translator (
		.clk                   (main_pll_sys_clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tristate_controller_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tristate_controller_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tristate_controller_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tristate_controller_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tristate_controller_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (tristate_controller_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (tristate_controller_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (tristate_controller_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (tristate_controller_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (tristate_controller_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (tristate_controller_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (85),
		.PKT_DATA_SIDEBAND_L       (85),
		.PKT_QOS_H                 (87),
		.PKT_QOS_L                 (87),
		.PKT_ADDR_SIDEBAND_H       (84),
		.PKT_ADDR_SIDEBAND_L       (84),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_data_master_translator_avalon_universal_master_0_agent (
		.clk              (main_pll_sys_clk_clk),                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (nios2_qsys_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (85),
		.PKT_DATA_SIDEBAND_L       (85),
		.PKT_QOS_H                 (87),
		.PKT_QOS_L                 (87),
		.PKT_ADDR_SIDEBAND_H       (84),
		.PKT_ADDR_SIDEBAND_L       (84),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (31),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (main_pll_sys_clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                                 //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                  //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                               //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                           //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                  //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (61),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (40),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (54),
		.PKT_BURST_SIZE_L          (52),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (70),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (63),
		.PKT_BURST_SIZE_L          (61),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                           //                .channel
		.rf_sink_ready           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                               //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                               //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                             //                .channel
		.rf_sink_ready           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) green_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                  //                .channel
		.rf_sink_ready           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_005_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_005_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_005_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_005_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_005_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_005_source0_channel),                                                      //                .channel
		.rf_sink_ready           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (70),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (63),
		.PKT_BURST_SIZE_L          (61),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_006_source0_ready),                                               //              cp.ready
		.cp_valid                (burst_adapter_006_source0_valid),                                               //                .valid
		.cp_data                 (burst_adapter_006_source0_data),                                                //                .data
		.cp_startofpacket        (burst_adapter_006_source0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_006_source0_endofpacket),                                         //                .endofpacket
		.cp_channel              (burst_adapter_006_source0_channel),                                             //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_007_source0_ready),                                                //              cp.ready
		.cp_valid                (burst_adapter_007_source0_valid),                                                //                .valid
		.cp_data                 (burst_adapter_007_source0_data),                                                 //                .data
		.cp_startofpacket        (burst_adapter_007_source0_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (burst_adapter_007_source0_endofpacket),                                          //                .endofpacket
		.cp_channel              (burst_adapter_007_source0_channel),                                              //                .channel
		.rf_sink_ready           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_008_source0_ready),                                               //              cp.ready
		.cp_valid                (burst_adapter_008_source0_valid),                                               //                .valid
		.cp_data                 (burst_adapter_008_source0_data),                                                //                .data
		.cp_startofpacket        (burst_adapter_008_source0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_008_source0_endofpacket),                                         //                .endofpacket
		.cp_channel              (burst_adapter_008_source0_channel),                                             //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_009_source0_ready),                                                                  //              cp.ready
		.cp_valid                (burst_adapter_009_source0_valid),                                                                  //                .valid
		.cp_data                 (burst_adapter_009_source0_data),                                                                   //                .data
		.cp_startofpacket        (burst_adapter_009_source0_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_009_source0_endofpacket),                                                            //                .endofpacket
		.cp_channel              (burst_adapter_009_source0_channel),                                                                //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) add_button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (add_button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (add_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (add_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (add_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (add_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (add_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (add_button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (add_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (add_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (add_button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (add_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (add_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (add_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (add_button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (add_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_010_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_010_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_010_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_010_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_010_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_010_source0_channel),                                                  //                .channel
		.rf_sink_ready           (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (add_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (add_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (add_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) remove_button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (remove_button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_011_source0_ready),                                                       //              cp.ready
		.cp_valid                (burst_adapter_011_source0_valid),                                                       //                .valid
		.cp_data                 (burst_adapter_011_source0_data),                                                        //                .data
		.cp_startofpacket        (burst_adapter_011_source0_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_011_source0_endofpacket),                                                 //                .endofpacket
		.cp_channel              (burst_adapter_011_source0_channel),                                                     //                .channel
		.rf_sink_ready           (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (remove_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (remove_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (remove_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cancel_button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cancel_button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_012_source0_ready),                                                       //              cp.ready
		.cp_valid                (burst_adapter_012_source0_valid),                                                       //                .valid
		.cp_data                 (burst_adapter_012_source0_data),                                                        //                .data
		.cp_startofpacket        (burst_adapter_012_source0_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_012_source0_endofpacket),                                                 //                .endofpacket
		.cp_channel              (burst_adapter_012_source0_channel),                                                     //                .channel
		.rf_sink_ready           (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cancel_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cancel_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) red_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_013_source0_ready),                                                  //              cp.ready
		.cp_valid                (burst_adapter_013_source0_valid),                                                  //                .valid
		.cp_data                 (burst_adapter_013_source0_data),                                                   //                .data
		.cp_startofpacket        (burst_adapter_013_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_013_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (burst_adapter_013_source0_channel),                                                //                .channel
		.rf_sink_ready           (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_014_source0_ready),                                                                           //              cp.ready
		.cp_valid                (burst_adapter_014_source0_valid),                                                                           //                .valid
		.cp_data                 (burst_adapter_014_source0_data),                                                                            //                .data
		.cp_startofpacket        (burst_adapter_014_source0_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_014_source0_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (burst_adapter_014_source0_channel),                                                                         //                .channel
		.rf_sink_ready           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_audio_clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_015_source0_ready),                                                                    //              cp.ready
		.cp_valid                (burst_adapter_015_source0_valid),                                                                    //                .valid
		.cp_data                 (burst_adapter_015_source0_data),                                                                     //                .data
		.cp_startofpacket        (burst_adapter_015_source0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_015_source0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (burst_adapter_015_source0_channel),                                                                  //                .channel
		.rf_sink_ready           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_audio_clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (main_pll_audio_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                                         // (terminated)
		.out_startofpacket (),                                                                                             // (terminated)
		.out_endofpacket   (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_016_source0_ready),                                                                          //              cp.ready
		.cp_valid                (burst_adapter_016_source0_valid),                                                                          //                .valid
		.cp_data                 (burst_adapter_016_source0_data),                                                                           //                .data
		.cp_startofpacket        (burst_adapter_016_source0_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (burst_adapter_016_source0_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (burst_adapter_016_source0_channel),                                                                        //                .channel
		.rf_sink_ready           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (88),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_017_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_017_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_017_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_017_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_017_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_017_source0_channel),                                                           //                .channel
		.rf_sink_ready           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (61),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (40),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (54),
		.PKT_BURST_SIZE_L          (52),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tristate_controller_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (main_pll_sys_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tristate_controller_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_018_source0_ready),                                                              //              cp.ready
		.cp_valid                (burst_adapter_018_source0_valid),                                                              //                .valid
		.cp_data                 (burst_adapter_018_source0_data),                                                               //                .data
		.cp_startofpacket        (burst_adapter_018_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (burst_adapter_018_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (burst_adapter_018_source0_channel),                                                            //                .channel
		.rf_sink_ready           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (main_pll_sys_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	niosII_system_addr_router addr_router (
		.sink_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	niosII_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                 //          .valid
		.src_data           (addr_router_001_src_data),                                                                  //          .data
		.src_channel        (addr_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	niosII_system_id_router id_router (
		.sink_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	niosII_system_id_router_001 id_router_001 (
		.sink_ready         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	niosII_system_id_router_002 id_router_002 (
		.sink_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	niosII_system_id_router_003 id_router_003 (
		.sink_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                                             //          .valid
		.src_data           (id_router_003_src_data),                                                              //          .data
		.src_channel        (id_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	niosII_system_id_router_003 id_router_004 (
		.sink_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                             //          .endofpacket
	);

	niosII_system_id_router id_router_005 (
		.sink_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                 //          .endofpacket
	);

	niosII_system_id_router_002 id_router_006 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                             //       src.ready
		.src_valid          (id_router_006_src_valid),                                             //          .valid
		.src_data           (id_router_006_src_data),                                              //          .data
		.src_channel        (id_router_006_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                        //          .endofpacket
	);

	niosII_system_id_router_003 id_router_007 (
		.sink_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                              //       src.ready
		.src_valid          (id_router_007_src_valid),                                              //          .valid
		.src_data           (id_router_007_src_data),                                               //          .data
		.src_channel        (id_router_007_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                         //          .endofpacket
	);

	niosII_system_id_router_003 id_router_008 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                             //       src.ready
		.src_valid          (id_router_008_src_valid),                                             //          .valid
		.src_data           (id_router_008_src_data),                                              //          .data
		.src_channel        (id_router_008_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                        //          .endofpacket
	);

	niosII_system_id_router_003 id_router_009 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                //          .valid
		.src_data           (id_router_009_src_data),                                                                 //          .data
		.src_channel        (id_router_009_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                           //          .endofpacket
	);

	niosII_system_id_router_003 id_router_010 (
		.sink_ready         (add_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (add_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (add_button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (add_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (add_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                  //       src.ready
		.src_valid          (id_router_010_src_valid),                                                  //          .valid
		.src_data           (id_router_010_src_data),                                                   //          .data
		.src_channel        (id_router_010_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                             //          .endofpacket
	);

	niosII_system_id_router_003 id_router_011 (
		.sink_ready         (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (remove_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                     //       src.ready
		.src_valid          (id_router_011_src_valid),                                                     //          .valid
		.src_data           (id_router_011_src_data),                                                      //          .data
		.src_channel        (id_router_011_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                //          .endofpacket
	);

	niosII_system_id_router_003 id_router_012 (
		.sink_ready         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cancel_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                     //       src.ready
		.src_valid          (id_router_012_src_valid),                                                     //          .valid
		.src_data           (id_router_012_src_data),                                                      //          .data
		.src_channel        (id_router_012_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                //          .endofpacket
	);

	niosII_system_id_router_003 id_router_013 (
		.sink_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                //       src.ready
		.src_valid          (id_router_013_src_valid),                                                //          .valid
		.src_data           (id_router_013_src_data),                                                 //          .data
		.src_channel        (id_router_013_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                           //          .endofpacket
	);

	niosII_system_id_router_003 id_router_014 (
		.sink_ready         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (barcode_scanner_ps2_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                         //          .valid
		.src_data           (id_router_014_src_data),                                                                          //          .data
		.src_channel        (id_router_014_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                                    //          .endofpacket
	);

	niosII_system_id_router_003 id_router_015 (
		.sink_ready         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_core_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_audio_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_015_src_valid),                                                                  //          .valid
		.src_data           (id_router_015_src_data),                                                                   //          .data
		.src_channel        (id_router_015_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_id_router_003 id_router_016 (
		.sink_ready         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_016_src_valid),                                                                        //          .valid
		.src_data           (id_router_016_src_data),                                                                         //          .data
		.src_channel        (id_router_016_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                                   //          .endofpacket
	);

	niosII_system_id_router_003 id_router_017 (
		.sink_ready         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dm9000a_if_ethernet_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                           //       src.ready
		.src_valid          (id_router_017_src_valid),                                                           //          .valid
		.src_data           (id_router_017_src_data),                                                            //          .data
		.src_channel        (id_router_017_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                      //          .endofpacket
	);

	niosII_system_id_router_018 id_router_018 (
		.sink_ready         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tristate_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (main_pll_sys_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                            //       src.ready
		.src_valid          (id_router_018_src_valid),                                                            //          .valid
		.src_data           (id_router_018_src_data),                                                             //          .data
		.src_channel        (id_router_018_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (main_pll_sys_clk_clk),           //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (main_pll_sys_clk_clk),               //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter (
		.clk                   (main_pll_sys_clk_clk),                //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_src_ready),              //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (40),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (54),
		.PKT_BURST_SIZE_L          (52),
		.PKT_BURST_TYPE_H          (56),
		.PKT_BURST_TYPE_L          (55),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (46),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (40),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_001 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),                 //     sink0.valid
		.sink0_data            (width_adapter_src_data),                  //          .data
		.sink0_channel         (width_adapter_src_channel),               //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),         //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),           //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),                 //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (63),
		.PKT_BURST_SIZE_L          (61),
		.PKT_BURST_TYPE_H          (65),
		.PKT_BURST_TYPE_L          (64),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (55),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (60),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter_002 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_003 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src3_valid),               //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src3_data),                //          .data
		.sink0_channel         (cmd_xbar_demux_src3_channel),             //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src3_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src3_endofpacket),         //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src3_ready),               //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_004 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src4_valid),               //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src4_data),                //          .data
		.sink0_channel         (cmd_xbar_demux_src4_channel),             //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src4_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src4_endofpacket),         //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src4_ready),               //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter_005 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_005_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_005_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_005_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_005_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_005_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_005_src_ready),              //          .ready
		.source0_valid         (burst_adapter_005_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_005_source0_data),          //          .data
		.source0_channel       (burst_adapter_005_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_005_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_005_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_005_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (63),
		.PKT_BURST_SIZE_L          (61),
		.PKT_BURST_TYPE_H          (65),
		.PKT_BURST_TYPE_L          (64),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (55),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (60),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter_006 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_006_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_006_source0_data),          //          .data
		.source0_channel       (burst_adapter_006_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_006_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_006_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_006_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_007 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src7_valid),               //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src7_data),                //          .data
		.sink0_channel         (cmd_xbar_demux_src7_channel),             //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src7_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src7_endofpacket),         //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src7_ready),               //          .ready
		.source0_valid         (burst_adapter_007_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_007_source0_data),          //          .data
		.source0_channel       (burst_adapter_007_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_007_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_007_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_007_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_008 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src8_valid),               //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src8_data),                //          .data
		.sink0_channel         (cmd_xbar_demux_src8_channel),             //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src8_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src8_endofpacket),         //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src8_ready),               //          .ready
		.source0_valid         (burst_adapter_008_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_008_source0_data),          //          .data
		.source0_channel       (burst_adapter_008_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_008_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_008_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_008_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_009 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src9_valid),               //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src9_data),                //          .data
		.sink0_channel         (cmd_xbar_demux_src9_channel),             //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src9_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src9_endofpacket),         //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src9_ready),               //          .ready
		.source0_valid         (burst_adapter_009_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_009_source0_data),          //          .data
		.source0_channel       (burst_adapter_009_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_009_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_009_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_009_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_010 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src10_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src10_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src10_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src10_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src10_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src10_ready),              //          .ready
		.source0_valid         (burst_adapter_010_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_010_source0_data),          //          .data
		.source0_channel       (burst_adapter_010_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_010_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_010_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_010_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_011 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src11_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src11_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src11_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src11_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src11_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src11_ready),              //          .ready
		.source0_valid         (burst_adapter_011_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_011_source0_data),          //          .data
		.source0_channel       (burst_adapter_011_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_011_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_011_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_011_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_012 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src12_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src12_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src12_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src12_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src12_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src12_ready),              //          .ready
		.source0_valid         (burst_adapter_012_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_012_source0_data),          //          .data
		.source0_channel       (burst_adapter_012_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_012_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_012_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_012_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_013 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src13_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src13_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src13_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src13_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src13_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src13_ready),              //          .ready
		.source0_valid         (burst_adapter_013_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_013_source0_data),          //          .data
		.source0_channel       (burst_adapter_013_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_013_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_013_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_013_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_014 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src14_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src14_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src14_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src14_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src14_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src14_ready),              //          .ready
		.source0_valid         (burst_adapter_014_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_014_source0_data),          //          .data
		.source0_channel       (burst_adapter_014_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_014_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_014_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_014_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_015 (
		.clk                   (main_pll_audio_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (crosser_out_valid),                       //     sink0.valid
		.sink0_data            (crosser_out_data),                        //          .data
		.sink0_channel         (crosser_out_channel),                     //          .channel
		.sink0_startofpacket   (crosser_out_startofpacket),               //          .startofpacket
		.sink0_endofpacket     (crosser_out_endofpacket),                 //          .endofpacket
		.sink0_ready           (crosser_out_ready),                       //          .ready
		.source0_valid         (burst_adapter_015_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_015_source0_data),          //          .data
		.source0_channel       (burst_adapter_015_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_015_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_015_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_015_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_016 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src16_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src16_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src16_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src16_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src16_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src16_ready),              //          .ready
		.source0_valid         (burst_adapter_016_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_016_source0_data),          //          .data
		.source0_channel       (burst_adapter_016_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_016_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_016_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_016_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (86),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (81),
		.PKT_BURST_SIZE_L          (79),
		.PKT_BURST_TYPE_H          (83),
		.PKT_BURST_TYPE_L          (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (73),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (69),
		.OUT_BURSTWRAP_H           (78),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter_017 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_src17_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_demux_src17_data),               //          .data
		.sink0_channel         (cmd_xbar_demux_src17_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_src17_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_src17_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_src17_ready),              //          .ready
		.source0_valid         (burst_adapter_017_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_017_source0_data),          //          .data
		.source0_channel       (burst_adapter_017_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_017_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_017_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_017_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (40),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (54),
		.PKT_BURST_SIZE_L          (52),
		.PKT_BURST_TYPE_H          (56),
		.PKT_BURST_TYPE_L          (55),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (46),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (40),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (31),
		.BURSTWRAP_CONST_VALUE     (31)
	) burst_adapter_018 (
		.clk                   (main_pll_sys_clk_clk),                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_006_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_006_src_data),              //          .data
		.sink0_channel         (width_adapter_006_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_006_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_006_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_006_src_ready),             //          .ready
		.source0_valid         (burst_adapter_018_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_018_source0_data),          //          .data
		.source0_channel       (burst_adapter_018_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_018_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_018_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_018_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (4),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                           // reset_in0.reset
		.reset_in1  (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~main_pll_sys_clk_reset_reset),            // reset_in2.reset
		.reset_in3  (~clock_27mhz_clk_in_reset_reset_n),        // reset_in3.reset
		.clk        (main_pll_sys_clk_clk),                     //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_in4  (1'b0),                                     // (terminated)
		.reset_in5  (1'b0),                                     // (terminated)
		.reset_in6  (1'b0),                                     // (terminated)
		.reset_in7  (1'b0),                                     // (terminated)
		.reset_in8  (1'b0),                                     // (terminated)
		.reset_in9  (1'b0),                                     // (terminated)
		.reset_in10 (1'b0),                                     // (terminated)
		.reset_in11 (1'b0),                                     // (terminated)
		.reset_in12 (1'b0),                                     // (terminated)
		.reset_in13 (1'b0),                                     // (terminated)
		.reset_in14 (1'b0),                                     // (terminated)
		.reset_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (4),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                           // reset_in0.reset
		.reset_in1  (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~main_pll_sys_clk_reset_reset),            // reset_in2.reset
		.reset_in3  (~clock_27mhz_clk_in_reset_reset_n),        // reset_in3.reset
		.clk        (main_pll_audio_clk_clk),                   //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),       // reset_out.reset
		.reset_in4  (1'b0),                                     // (terminated)
		.reset_in5  (1'b0),                                     // (terminated)
		.reset_in6  (1'b0),                                     // (terminated)
		.reset_in7  (1'b0),                                     // (terminated)
		.reset_in8  (1'b0),                                     // (terminated)
		.reset_in9  (1'b0),                                     // (terminated)
		.reset_in10 (1'b0),                                     // (terminated)
		.reset_in11 (1'b0),                                     // (terminated)
		.reset_in12 (1'b0),                                     // (terminated)
		.reset_in13 (1'b0),                                     // (terminated)
		.reset_in14 (1'b0),                                     // (terminated)
		.reset_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (4),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                           // reset_in0.reset
		.reset_in1  (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~main_pll_sys_clk_reset_reset),            // reset_in2.reset
		.reset_in3  (~clock_27mhz_clk_in_reset_reset_n),        // reset_in3.reset
		.clk        (clk_clk),                                  //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),       // reset_out.reset
		.reset_in4  (1'b0),                                     // (terminated)
		.reset_in5  (1'b0),                                     // (terminated)
		.reset_in6  (1'b0),                                     // (terminated)
		.reset_in7  (1'b0),                                     // (terminated)
		.reset_in8  (1'b0),                                     // (terminated)
		.reset_in9  (1'b0),                                     // (terminated)
		.reset_in10 (1'b0),                                     // (terminated)
		.reset_in11 (1'b0),                                     // (terminated)
		.reset_in12 (1'b0),                                     // (terminated)
		.reset_in13 (1'b0),                                     // (terminated)
		.reset_in14 (1'b0),                                     // (terminated)
		.reset_in15 (1'b0)                                      // (terminated)
	);

	niosII_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (main_pll_sys_clk_clk),               //        clk.clk
		.reset               (rst_controller_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_cmd_src_channel),            //           .channel
		.sink_data           (limiter_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_src18_endofpacket)    //           .endofpacket
	);

	niosII_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (main_pll_sys_clk_clk),                  //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //           .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_018 (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_018_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_018_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_018_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_018_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_018_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_018_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src18_ready),            //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src18_valid),            //          .valid
		.sink0_channel       (cmd_xbar_demux_src18_channel),          //          .channel
		.sink0_data          (cmd_xbar_demux_src18_data),             //          .data
		.sink0_startofpacket (cmd_xbar_demux_src18_startofpacket),    //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src18_endofpacket),      //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (main_pll_sys_clk_clk),              //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_003 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_004 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_007 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_008 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_009 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_010 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_011 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_012 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_013 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_014 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_015 (
		.clk                (main_pll_audio_clk_clk),                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_016 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_001 rsp_xbar_demux_017 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_018 (
		.clk                (main_pll_sys_clk_clk),                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_007_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_007_src_channel),         //          .channel
		.sink_data          (width_adapter_007_src_data),            //          .data
		.sink_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_007_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_018_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (main_pll_sys_clk_clk),                  //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (crosser_001_out_ready),                 //    sink15.ready
		.sink15_valid         (crosser_001_out_valid),                 //          .valid
		.sink15_channel       (crosser_001_out_channel),               //          .channel
		.sink15_data          (crosser_001_out_data),                  //          .data
		.sink15_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink15_endofpacket   (crosser_001_out_endofpacket),           //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (main_pll_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_002_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_005_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_006_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_018_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (81),
		.IN_PKT_BURST_SIZE_L           (79),
		.IN_PKT_RESPONSE_STATUS_H      (107),
		.IN_PKT_RESPONSE_STATUS_L      (106),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (83),
		.IN_PKT_BURST_TYPE_L           (82),
		.IN_ST_DATA_W                  (108),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (45),
		.OUT_PKT_BYTE_CNT_L            (40),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_PKT_BURST_SIZE_H          (54),
		.OUT_PKT_BURST_SIZE_L          (52),
		.OUT_PKT_RESPONSE_STATUS_H     (80),
		.OUT_PKT_RESPONSE_STATUS_L     (79),
		.OUT_PKT_TRANS_EXCLUSIVE       (39),
		.OUT_PKT_BURST_TYPE_H          (56),
		.OUT_PKT_BURST_TYPE_L          (55),
		.OUT_ST_DATA_W                 (81),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (main_pll_sys_clk_clk),              //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src1_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (45),
		.IN_PKT_BYTE_CNT_L             (40),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (46),
		.IN_PKT_BURST_SIZE_H           (54),
		.IN_PKT_BURST_SIZE_L           (52),
		.IN_PKT_RESPONSE_STATUS_H      (80),
		.IN_PKT_RESPONSE_STATUS_L      (79),
		.IN_PKT_TRANS_EXCLUSIVE        (39),
		.IN_PKT_BURST_TYPE_H           (56),
		.IN_PKT_BURST_TYPE_L           (55),
		.IN_ST_DATA_W                  (81),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (81),
		.OUT_PKT_BURST_SIZE_L          (79),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (83),
		.OUT_PKT_BURST_TYPE_L          (82),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_001 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (81),
		.IN_PKT_BURST_SIZE_L           (79),
		.IN_PKT_RESPONSE_STATUS_H      (107),
		.IN_PKT_RESPONSE_STATUS_L      (106),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (83),
		.IN_PKT_BURST_TYPE_L           (82),
		.IN_ST_DATA_W                  (108),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (54),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (63),
		.OUT_PKT_BURST_SIZE_L          (61),
		.OUT_PKT_RESPONSE_STATUS_H     (89),
		.OUT_PKT_RESPONSE_STATUS_L     (88),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (65),
		.OUT_PKT_BURST_TYPE_L          (64),
		.OUT_ST_DATA_W                 (90),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (54),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (60),
		.IN_PKT_BURSTWRAP_L            (55),
		.IN_PKT_BURST_SIZE_H           (63),
		.IN_PKT_BURST_SIZE_L           (61),
		.IN_PKT_RESPONSE_STATUS_H      (89),
		.IN_PKT_RESPONSE_STATUS_L      (88),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (65),
		.IN_PKT_BURST_TYPE_L           (64),
		.IN_ST_DATA_W                  (90),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (81),
		.OUT_PKT_BURST_SIZE_L          (79),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (83),
		.OUT_PKT_BURST_TYPE_L          (82),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_003 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (81),
		.IN_PKT_BURST_SIZE_L           (79),
		.IN_PKT_RESPONSE_STATUS_H      (107),
		.IN_PKT_RESPONSE_STATUS_L      (106),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (83),
		.IN_PKT_BURST_TYPE_L           (82),
		.IN_ST_DATA_W                  (108),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (54),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (63),
		.OUT_PKT_BURST_SIZE_L          (61),
		.OUT_PKT_RESPONSE_STATUS_H     (89),
		.OUT_PKT_RESPONSE_STATUS_L     (88),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (65),
		.OUT_PKT_BURST_TYPE_L          (64),
		.OUT_ST_DATA_W                 (90),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_006_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_006_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_006_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_006_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_006_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_006_src_data),           //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_004_src_data),          //          .data
		.out_channel          (width_adapter_004_src_channel),       //          .channel
		.out_valid            (width_adapter_004_src_valid),         //          .valid
		.out_ready            (width_adapter_004_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (54),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (60),
		.IN_PKT_BURSTWRAP_L            (55),
		.IN_PKT_BURST_SIZE_H           (63),
		.IN_PKT_BURST_SIZE_L           (61),
		.IN_PKT_RESPONSE_STATUS_H      (89),
		.IN_PKT_RESPONSE_STATUS_L      (88),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (65),
		.IN_PKT_BURST_TYPE_L           (64),
		.IN_ST_DATA_W                  (90),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (81),
		.OUT_PKT_BURST_SIZE_L          (79),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (83),
		.OUT_PKT_BURST_TYPE_L          (82),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_005 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_006_src_valid),             //      sink.valid
		.in_channel           (id_router_006_src_channel),           //          .channel
		.in_startofpacket     (id_router_006_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_006_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_006_src_ready),             //          .ready
		.in_data              (id_router_006_src_data),              //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_005_src_data),          //          .data
		.out_channel          (width_adapter_005_src_channel),       //          .channel
		.out_valid            (width_adapter_005_src_valid),         //          .valid
		.out_ready            (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (72),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (73),
		.IN_PKT_BURST_SIZE_H           (81),
		.IN_PKT_BURST_SIZE_L           (79),
		.IN_PKT_RESPONSE_STATUS_H      (107),
		.IN_PKT_RESPONSE_STATUS_L      (106),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (83),
		.IN_PKT_BURST_TYPE_L           (82),
		.IN_ST_DATA_W                  (108),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (45),
		.OUT_PKT_BYTE_CNT_L            (40),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_PKT_BURST_SIZE_H          (54),
		.OUT_PKT_BURST_SIZE_L          (52),
		.OUT_PKT_RESPONSE_STATUS_H     (80),
		.OUT_PKT_RESPONSE_STATUS_L     (79),
		.OUT_PKT_TRANS_EXCLUSIVE       (39),
		.OUT_PKT_BURST_TYPE_H          (56),
		.OUT_PKT_BURST_TYPE_L          (55),
		.OUT_ST_DATA_W                 (81),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_006 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_018_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_018_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_018_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_018_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_018_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_018_src_data),           //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_006_src_data),          //          .data
		.out_channel          (width_adapter_006_src_channel),       //          .channel
		.out_valid            (width_adapter_006_src_valid),         //          .valid
		.out_ready            (width_adapter_006_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (45),
		.IN_PKT_BYTE_CNT_L             (40),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (46),
		.IN_PKT_BURST_SIZE_H           (54),
		.IN_PKT_BURST_SIZE_L           (52),
		.IN_PKT_RESPONSE_STATUS_H      (80),
		.IN_PKT_RESPONSE_STATUS_L      (79),
		.IN_PKT_TRANS_EXCLUSIVE        (39),
		.IN_PKT_BURST_TYPE_H           (56),
		.IN_PKT_BURST_TYPE_L           (55),
		.IN_ST_DATA_W                  (81),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (72),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (81),
		.OUT_PKT_BURST_SIZE_L          (79),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (83),
		.OUT_PKT_BURST_TYPE_L          (82),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_007 (
		.clk                  (main_pll_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_018_src_valid),             //      sink.valid
		.in_channel           (id_router_018_src_channel),           //          .channel
		.in_startofpacket     (id_router_018_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_018_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_018_src_ready),             //          .ready
		.in_data              (id_router_018_src_data),              //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_007_src_data),          //          .data
		.out_channel          (width_adapter_007_src_channel),       //          .channel
		.out_valid            (width_adapter_007_src_valid),         //          .valid
		.out_ready            (width_adapter_007_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (108),
		.BITS_PER_SYMBOL     (108),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (main_pll_sys_clk_clk),               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (main_pll_audio_clk_clk),             //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src15_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_src15_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_src15_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src15_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_src15_channel),       //              .channel
		.in_data           (cmd_xbar_demux_src15_data),          //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (108),
		.BITS_PER_SYMBOL     (108),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (19),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (main_pll_audio_clk_clk),                //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (main_pll_sys_clk_clk),                  //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_015_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_015_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_015_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_015_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	niosII_system_irq_mapper irq_mapper (
		.clk           (main_pll_sys_clk_clk),           //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (main_pll_audio_clk_clk),             //       receiver_clk.clk
		.sender_clk     (main_pll_sys_clk_clk),               //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

endmodule
